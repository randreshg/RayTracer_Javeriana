-- megafunction wizard: %ALTFP_ADD_SUB%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_add_sub 

-- ============================================================
-- File Name: addSub.vhd
-- Megafunction Name(s):
-- 			altfp_add_sub
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_add_sub CBX_AUTO_BLACKBOX="ALL" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone IV E" DIRECTION="VARIABLE" OPTIMIZE="SPEED" PIPELINE=7 REDUCED_FUNCTIONALITY="NO" WIDTH_EXP=8 WIDTH_MAN=23 add_sub clock dataa datab result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_altfp_add_sub 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=1 SHIFTDIR="LEFT" WIDTH=26 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = reg 27 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altbarrel_shift_35e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END addSub_altbarrel_shift_35e;

 ARCHITECTURE RTL OF addSub_altbarrel_shift_35e IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w695w696w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w691w692w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w716w717w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w712w713w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w738w739w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w734w735w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w760w761w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w756w757w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w782w783w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w778w779w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w687w688w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w708w709w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w730w731w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w752w753w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w774w775w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range682w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range682w691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range703w716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range703w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range725w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range725w734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range747w760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range747w756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range769w782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range769w778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_dir_w_range679w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_dir_w_range701w715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_dir_w_range722w737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_dir_w_range744w759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_dir_w_range766w781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range682w687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range703w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range725w730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range747w752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_sel_w_range769w774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range682w695w696w697w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range703w716w717w718w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range725w738w739w740w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range747w760w761w762w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range769w782w783w784w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w698w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w719w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w741w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w763w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w785w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (155 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (129 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w690w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w693w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w711w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w714w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w733w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w736w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w755w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w758w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w777w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w780w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_dir_w_range679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_dir_w_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_dir_w_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_dir_w_range744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_dir_w_range766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sbit_w_range742w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sbit_w_range764w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sbit_w_range677w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sbit_w_range700w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sbit_w_range720w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sel_w_range682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sel_w_range703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sel_w_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sel_w_range747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_sel_w_range769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lbarrel_shift_w_smux_w_range773w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w695w696w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range682w695w(0) AND wire_lbarrel_shift_w693w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w691w692w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range682w691w(0) AND wire_lbarrel_shift_w690w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w716w717w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range703w716w(0) AND wire_lbarrel_shift_w714w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w712w713w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range703w712w(0) AND wire_lbarrel_shift_w711w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w738w739w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range725w738w(0) AND wire_lbarrel_shift_w736w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w734w735w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range725w734w(0) AND wire_lbarrel_shift_w733w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w760w761w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range747w760w(0) AND wire_lbarrel_shift_w758w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w756w757w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range747w756w(0) AND wire_lbarrel_shift_w755w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w782w783w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range769w782w(0) AND wire_lbarrel_shift_w780w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w778w779w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range769w778w(0) AND wire_lbarrel_shift_w777w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w687w688w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range682w687w(0) AND wire_lbarrel_shift_w_sbit_w_range677w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w708w709w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range703w708w(0) AND wire_lbarrel_shift_w_sbit_w_range700w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w730w731w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range725w730w(0) AND wire_lbarrel_shift_w_sbit_w_range720w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w752w753w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range747w752w(0) AND wire_lbarrel_shift_w_sbit_w_range742w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w774w775w(i) <= wire_lbarrel_shift_w_lg_w_sel_w_range769w774w(0) AND wire_lbarrel_shift_w_sbit_w_range764w(i);
	END GENERATE loop14;
	wire_lbarrel_shift_w_lg_w_sel_w_range682w695w(0) <= wire_lbarrel_shift_w_sel_w_range682w(0) AND wire_lbarrel_shift_w_lg_w_dir_w_range679w694w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range682w691w(0) <= wire_lbarrel_shift_w_sel_w_range682w(0) AND wire_lbarrel_shift_w_dir_w_range679w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range703w716w(0) <= wire_lbarrel_shift_w_sel_w_range703w(0) AND wire_lbarrel_shift_w_lg_w_dir_w_range701w715w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range703w712w(0) <= wire_lbarrel_shift_w_sel_w_range703w(0) AND wire_lbarrel_shift_w_dir_w_range701w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range725w738w(0) <= wire_lbarrel_shift_w_sel_w_range725w(0) AND wire_lbarrel_shift_w_lg_w_dir_w_range722w737w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range725w734w(0) <= wire_lbarrel_shift_w_sel_w_range725w(0) AND wire_lbarrel_shift_w_dir_w_range722w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range747w760w(0) <= wire_lbarrel_shift_w_sel_w_range747w(0) AND wire_lbarrel_shift_w_lg_w_dir_w_range744w759w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range747w756w(0) <= wire_lbarrel_shift_w_sel_w_range747w(0) AND wire_lbarrel_shift_w_dir_w_range744w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range769w782w(0) <= wire_lbarrel_shift_w_sel_w_range769w(0) AND wire_lbarrel_shift_w_lg_w_dir_w_range766w781w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range769w778w(0) <= wire_lbarrel_shift_w_sel_w_range769w(0) AND wire_lbarrel_shift_w_dir_w_range766w(0);
	wire_lbarrel_shift_w_lg_w_dir_w_range679w694w(0) <= NOT wire_lbarrel_shift_w_dir_w_range679w(0);
	wire_lbarrel_shift_w_lg_w_dir_w_range701w715w(0) <= NOT wire_lbarrel_shift_w_dir_w_range701w(0);
	wire_lbarrel_shift_w_lg_w_dir_w_range722w737w(0) <= NOT wire_lbarrel_shift_w_dir_w_range722w(0);
	wire_lbarrel_shift_w_lg_w_dir_w_range744w759w(0) <= NOT wire_lbarrel_shift_w_dir_w_range744w(0);
	wire_lbarrel_shift_w_lg_w_dir_w_range766w781w(0) <= NOT wire_lbarrel_shift_w_dir_w_range766w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range682w687w(0) <= NOT wire_lbarrel_shift_w_sel_w_range682w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range703w708w(0) <= NOT wire_lbarrel_shift_w_sel_w_range703w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range725w730w(0) <= NOT wire_lbarrel_shift_w_sel_w_range725w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range747w752w(0) <= NOT wire_lbarrel_shift_w_sel_w_range747w(0);
	wire_lbarrel_shift_w_lg_w_sel_w_range769w774w(0) <= NOT wire_lbarrel_shift_w_sel_w_range769w(0);
	loop15 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range682w695w696w697w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w695w696w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w691w692w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range703w716w717w718w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w716w717w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w712w713w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range725w738w739w740w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w738w739w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w734w735w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range747w760w761w762w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w760w761w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w756w757w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range769w782w783w784w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w782w783w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w778w779w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w698w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range682w695w696w697w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range682w687w688w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w719w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range703w716w717w718w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range703w708w709w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w741w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range725w738w739w740w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range725w730w731w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w763w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range747w760w761w762w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range747w752w753w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 25 GENERATE 
		wire_lbarrel_shift_w785w(i) <= wire_lbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range769w782w783w784w(i) OR wire_lbarrel_shift_w_lg_w_lg_w_sel_w_range769w774w775w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(0) & dir_w(3 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(155 DOWNTO 130);
	sbit_w <= ( sbit_piper1d & smux_w(103 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_lbarrel_shift_w785w & wire_lbarrel_shift_w763w & wire_lbarrel_shift_w741w & wire_lbarrel_shift_w719w & wire_lbarrel_shift_w698w);
	wire_lbarrel_shift_w690w <= ( pad_w(0) & sbit_w(25 DOWNTO 1));
	wire_lbarrel_shift_w693w <= ( sbit_w(24 DOWNTO 0) & pad_w(0));
	wire_lbarrel_shift_w711w <= ( pad_w(1 DOWNTO 0) & sbit_w(51 DOWNTO 28));
	wire_lbarrel_shift_w714w <= ( sbit_w(49 DOWNTO 26) & pad_w(1 DOWNTO 0));
	wire_lbarrel_shift_w733w <= ( pad_w(3 DOWNTO 0) & sbit_w(77 DOWNTO 56));
	wire_lbarrel_shift_w736w <= ( sbit_w(73 DOWNTO 52) & pad_w(3 DOWNTO 0));
	wire_lbarrel_shift_w755w <= ( pad_w(7 DOWNTO 0) & sbit_w(103 DOWNTO 86));
	wire_lbarrel_shift_w758w <= ( sbit_w(95 DOWNTO 78) & pad_w(7 DOWNTO 0));
	wire_lbarrel_shift_w777w <= ( pad_w(15 DOWNTO 0) & sbit_w(129 DOWNTO 120));
	wire_lbarrel_shift_w780w <= ( sbit_w(113 DOWNTO 104) & pad_w(15 DOWNTO 0));
	wire_lbarrel_shift_w_dir_w_range679w(0) <= dir_w(0);
	wire_lbarrel_shift_w_dir_w_range701w(0) <= dir_w(1);
	wire_lbarrel_shift_w_dir_w_range722w(0) <= dir_w(2);
	wire_lbarrel_shift_w_dir_w_range744w(0) <= dir_w(3);
	wire_lbarrel_shift_w_dir_w_range766w(0) <= dir_w(4);
	wire_lbarrel_shift_w_sbit_w_range742w <= sbit_w(103 DOWNTO 78);
	wire_lbarrel_shift_w_sbit_w_range764w <= sbit_w(129 DOWNTO 104);
	wire_lbarrel_shift_w_sbit_w_range677w <= sbit_w(25 DOWNTO 0);
	wire_lbarrel_shift_w_sbit_w_range700w <= sbit_w(51 DOWNTO 26);
	wire_lbarrel_shift_w_sbit_w_range720w <= sbit_w(77 DOWNTO 52);
	wire_lbarrel_shift_w_sel_w_range682w(0) <= sel_w(0);
	wire_lbarrel_shift_w_sel_w_range703w(0) <= sel_w(1);
	wire_lbarrel_shift_w_sel_w_range725w(0) <= sel_w(2);
	wire_lbarrel_shift_w_sel_w_range747w(0) <= sel_w(3);
	wire_lbarrel_shift_w_sel_w_range769w(0) <= sel_w(4);
	wire_lbarrel_shift_w_smux_w_range773w <= smux_w(129 DOWNTO 104);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe(0) <= ( dir_w(4));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_lbarrel_shift_w_smux_w_range773w;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --addSub_altbarrel_shift_35e


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" SHIFTDIR="RIGHT" WIDTH=26 WIDTHDIST=5 data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altbarrel_shift_olb IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END addSub_altbarrel_shift_olb;

 ARCHITECTURE RTL OF addSub_altbarrel_shift_olb IS

	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w809w810w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w805w806w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w830w831w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w826w827w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w852w853w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w848w849w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w874w875w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w870w871w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w896w897w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w892w893w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w801w802w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w822w823w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w844w845w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w866w867w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w888w889w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range796w809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range796w805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range817w830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range817w826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range839w852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range839w848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range861w874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range861w870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range883w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range883w892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_dir_w_range793w808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_dir_w_range815w829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_dir_w_range836w851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_dir_w_range858w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_dir_w_range880w895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range796w801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range817w822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range839w844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range861w866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_sel_w_range883w888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range796w809w810w811w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range817w830w831w832w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range839w852w853w854w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range861w874w875w876w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range883w896w897w898w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w812w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w833w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w855w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w877w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w899w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (155 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (129 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w804w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w807w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w825w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w828w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w847w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w850w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w869w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w872w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w891w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w894w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_dir_w_range793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_dir_w_range815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_dir_w_range836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_dir_w_range858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_dir_w_range880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sbit_w_range856w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sbit_w_range878w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sbit_w_range791w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sbit_w_range814w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sbit_w_range834w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sel_w_range796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sel_w_range817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sel_w_range839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sel_w_range861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_w_sel_w_range883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	loop25 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w809w810w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range796w809w(0) AND wire_rbarrel_shift_w807w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w805w806w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range796w805w(0) AND wire_rbarrel_shift_w804w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w830w831w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range817w830w(0) AND wire_rbarrel_shift_w828w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w826w827w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range817w826w(0) AND wire_rbarrel_shift_w825w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w852w853w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range839w852w(0) AND wire_rbarrel_shift_w850w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w848w849w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range839w848w(0) AND wire_rbarrel_shift_w847w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w874w875w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range861w874w(0) AND wire_rbarrel_shift_w872w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w870w871w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range861w870w(0) AND wire_rbarrel_shift_w869w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w896w897w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range883w896w(0) AND wire_rbarrel_shift_w894w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w892w893w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range883w892w(0) AND wire_rbarrel_shift_w891w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w801w802w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range796w801w(0) AND wire_rbarrel_shift_w_sbit_w_range791w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w822w823w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range817w822w(0) AND wire_rbarrel_shift_w_sbit_w_range814w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w844w845w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range839w844w(0) AND wire_rbarrel_shift_w_sbit_w_range834w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w866w867w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range861w866w(0) AND wire_rbarrel_shift_w_sbit_w_range856w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w888w889w(i) <= wire_rbarrel_shift_w_lg_w_sel_w_range883w888w(0) AND wire_rbarrel_shift_w_sbit_w_range878w(i);
	END GENERATE loop39;
	wire_rbarrel_shift_w_lg_w_sel_w_range796w809w(0) <= wire_rbarrel_shift_w_sel_w_range796w(0) AND wire_rbarrel_shift_w_lg_w_dir_w_range793w808w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range796w805w(0) <= wire_rbarrel_shift_w_sel_w_range796w(0) AND wire_rbarrel_shift_w_dir_w_range793w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range817w830w(0) <= wire_rbarrel_shift_w_sel_w_range817w(0) AND wire_rbarrel_shift_w_lg_w_dir_w_range815w829w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range817w826w(0) <= wire_rbarrel_shift_w_sel_w_range817w(0) AND wire_rbarrel_shift_w_dir_w_range815w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range839w852w(0) <= wire_rbarrel_shift_w_sel_w_range839w(0) AND wire_rbarrel_shift_w_lg_w_dir_w_range836w851w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range839w848w(0) <= wire_rbarrel_shift_w_sel_w_range839w(0) AND wire_rbarrel_shift_w_dir_w_range836w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range861w874w(0) <= wire_rbarrel_shift_w_sel_w_range861w(0) AND wire_rbarrel_shift_w_lg_w_dir_w_range858w873w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range861w870w(0) <= wire_rbarrel_shift_w_sel_w_range861w(0) AND wire_rbarrel_shift_w_dir_w_range858w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range883w896w(0) <= wire_rbarrel_shift_w_sel_w_range883w(0) AND wire_rbarrel_shift_w_lg_w_dir_w_range880w895w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range883w892w(0) <= wire_rbarrel_shift_w_sel_w_range883w(0) AND wire_rbarrel_shift_w_dir_w_range880w(0);
	wire_rbarrel_shift_w_lg_w_dir_w_range793w808w(0) <= NOT wire_rbarrel_shift_w_dir_w_range793w(0);
	wire_rbarrel_shift_w_lg_w_dir_w_range815w829w(0) <= NOT wire_rbarrel_shift_w_dir_w_range815w(0);
	wire_rbarrel_shift_w_lg_w_dir_w_range836w851w(0) <= NOT wire_rbarrel_shift_w_dir_w_range836w(0);
	wire_rbarrel_shift_w_lg_w_dir_w_range858w873w(0) <= NOT wire_rbarrel_shift_w_dir_w_range858w(0);
	wire_rbarrel_shift_w_lg_w_dir_w_range880w895w(0) <= NOT wire_rbarrel_shift_w_dir_w_range880w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range796w801w(0) <= NOT wire_rbarrel_shift_w_sel_w_range796w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range817w822w(0) <= NOT wire_rbarrel_shift_w_sel_w_range817w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range839w844w(0) <= NOT wire_rbarrel_shift_w_sel_w_range839w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range861w866w(0) <= NOT wire_rbarrel_shift_w_sel_w_range861w(0);
	wire_rbarrel_shift_w_lg_w_sel_w_range883w888w(0) <= NOT wire_rbarrel_shift_w_sel_w_range883w(0);
	loop40 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range796w809w810w811w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w809w810w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w805w806w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range817w830w831w832w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w830w831w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w826w827w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range839w852w853w854w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w852w853w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w848w849w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range861w874w875w876w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w874w875w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w870w871w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range883w896w897w898w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w896w897w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w892w893w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w812w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range796w809w810w811w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range796w801w802w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w833w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range817w830w831w832w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range817w822w823w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w855w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range839w852w853w854w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range839w844w845w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w877w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range861w874w875w876w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range861w866w867w(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 25 GENERATE 
		wire_rbarrel_shift_w899w(i) <= wire_rbarrel_shift_w_lg_w_lg_w_lg_w_sel_w_range883w896w897w898w(i) OR wire_rbarrel_shift_w_lg_w_lg_w_sel_w_range883w888w889w(i);
	END GENERATE loop49;
	dir_w <= ( dir_w(4 DOWNTO 0) & direction_w);
	direction_w <= '1';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(155 DOWNTO 130);
	sbit_w <= ( smux_w(129 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_rbarrel_shift_w899w & wire_rbarrel_shift_w877w & wire_rbarrel_shift_w855w & wire_rbarrel_shift_w833w & wire_rbarrel_shift_w812w);
	wire_rbarrel_shift_w804w <= ( pad_w(0) & sbit_w(25 DOWNTO 1));
	wire_rbarrel_shift_w807w <= ( sbit_w(24 DOWNTO 0) & pad_w(0));
	wire_rbarrel_shift_w825w <= ( pad_w(1 DOWNTO 0) & sbit_w(51 DOWNTO 28));
	wire_rbarrel_shift_w828w <= ( sbit_w(49 DOWNTO 26) & pad_w(1 DOWNTO 0));
	wire_rbarrel_shift_w847w <= ( pad_w(3 DOWNTO 0) & sbit_w(77 DOWNTO 56));
	wire_rbarrel_shift_w850w <= ( sbit_w(73 DOWNTO 52) & pad_w(3 DOWNTO 0));
	wire_rbarrel_shift_w869w <= ( pad_w(7 DOWNTO 0) & sbit_w(103 DOWNTO 86));
	wire_rbarrel_shift_w872w <= ( sbit_w(95 DOWNTO 78) & pad_w(7 DOWNTO 0));
	wire_rbarrel_shift_w891w <= ( pad_w(15 DOWNTO 0) & sbit_w(129 DOWNTO 120));
	wire_rbarrel_shift_w894w <= ( sbit_w(113 DOWNTO 104) & pad_w(15 DOWNTO 0));
	wire_rbarrel_shift_w_dir_w_range793w(0) <= dir_w(0);
	wire_rbarrel_shift_w_dir_w_range815w(0) <= dir_w(1);
	wire_rbarrel_shift_w_dir_w_range836w(0) <= dir_w(2);
	wire_rbarrel_shift_w_dir_w_range858w(0) <= dir_w(3);
	wire_rbarrel_shift_w_dir_w_range880w(0) <= dir_w(4);
	wire_rbarrel_shift_w_sbit_w_range856w <= sbit_w(103 DOWNTO 78);
	wire_rbarrel_shift_w_sbit_w_range878w <= sbit_w(129 DOWNTO 104);
	wire_rbarrel_shift_w_sbit_w_range791w <= sbit_w(25 DOWNTO 0);
	wire_rbarrel_shift_w_sbit_w_range814w <= sbit_w(51 DOWNTO 26);
	wire_rbarrel_shift_w_sbit_w_range834w <= sbit_w(77 DOWNTO 52);
	wire_rbarrel_shift_w_sel_w_range796w(0) <= sel_w(0);
	wire_rbarrel_shift_w_sel_w_range817w(0) <= sel_w(1);
	wire_rbarrel_shift_w_sel_w_range839w(0) <= sel_w(2);
	wire_rbarrel_shift_w_sel_w_range861w(0) <= sel_w(3);
	wire_rbarrel_shift_w_sel_w_range883w(0) <= sel_w(4);

 END RTL; --addSub_altbarrel_shift_olb


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --addSub_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero934w935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero936w937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero934w & wire_altpriority_encoder14_w_lg_w_lg_zero936w937w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  addSub_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	wire_altpriority_encoder14_w_lg_w_lg_zero934w935w(0) <= wire_altpriority_encoder14_w_lg_zero934w(0) AND wire_altpriority_encoder14_q(0);
	wire_altpriority_encoder14_w_lg_zero936w(0) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(0);
	wire_altpriority_encoder14_w_lg_zero934w(0) <= NOT wire_altpriority_encoder14_zero;
	wire_altpriority_encoder14_w_lg_w_lg_zero936w937w(0) <= wire_altpriority_encoder14_w_lg_zero936w(0) OR wire_altpriority_encoder14_w_lg_w_lg_zero934w935w(0);
	altpriority_encoder14 :  addSub_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --addSub_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_be8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero924w925w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero926w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero926w927w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero924w & wire_altpriority_encoder12_w_lg_w_lg_zero926w927w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  addSub_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	loop50 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero924w925w(i) <= wire_altpriority_encoder12_w_lg_zero924w(0) AND wire_altpriority_encoder12_q(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder12_w_lg_zero926w(i) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(i);
	END GENERATE loop51;
	wire_altpriority_encoder12_w_lg_zero924w(0) <= NOT wire_altpriority_encoder12_zero;
	loop52 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero926w927w(i) <= wire_altpriority_encoder12_w_lg_zero926w(i) OR wire_altpriority_encoder12_w_lg_w_lg_zero924w925w(i);
	END GENERATE loop52;
	altpriority_encoder12 :  addSub_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --addSub_altpriority_encoder_be8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --addSub_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero959w960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero961w962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero959w & wire_altpriority_encoder18_w_lg_w_lg_zero961w962w);
	altpriority_encoder17 :  addSub_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	wire_altpriority_encoder18_w_lg_w_lg_zero959w960w(0) <= wire_altpriority_encoder18_w_lg_zero959w(0) AND wire_altpriority_encoder18_q(0);
	wire_altpriority_encoder18_w_lg_zero961w(0) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(0);
	wire_altpriority_encoder18_w_lg_zero959w(0) <= NOT wire_altpriority_encoder18_zero;
	wire_altpriority_encoder18_w_lg_w_lg_zero961w962w(0) <= wire_altpriority_encoder18_w_lg_zero961w(0) OR wire_altpriority_encoder18_w_lg_w_lg_zero959w960w(0);
	altpriority_encoder18 :  addSub_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --addSub_altpriority_encoder_6v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero950w951w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero952w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero952w953w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero950w & wire_altpriority_encoder16_w_lg_w_lg_zero952w953w);
	altpriority_encoder15 :  addSub_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder15_q
	  );
	loop53 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero950w951w(i) <= wire_altpriority_encoder16_w_lg_zero950w(0) AND wire_altpriority_encoder16_q(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_zero952w(i) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(i);
	END GENERATE loop54;
	wire_altpriority_encoder16_w_lg_zero950w(0) <= NOT wire_altpriority_encoder16_zero;
	loop55 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero952w953w(i) <= wire_altpriority_encoder16_w_lg_zero952w(i) OR wire_altpriority_encoder16_w_lg_w_lg_zero950w951w(i);
	END GENERATE loop55;
	altpriority_encoder16 :  addSub_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --addSub_altpriority_encoder_bv7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_r08;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero915w916w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero917w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero917w918w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 COMPONENT  addSub_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero915w & wire_altpriority_encoder10_w_lg_w_lg_zero917w918w);
	loop56 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero915w916w(i) <= wire_altpriority_encoder10_w_lg_zero915w(0) AND wire_altpriority_encoder10_q(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder10_w_lg_zero917w(i) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(i);
	END GENERATE loop57;
	wire_altpriority_encoder10_w_lg_zero915w(0) <= NOT wire_altpriority_encoder10_zero;
	loop58 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero917w918w(i) <= wire_altpriority_encoder10_w_lg_zero917w(i) OR wire_altpriority_encoder10_w_lg_w_lg_zero915w916w(i);
	END GENERATE loop58;
	altpriority_encoder10 :  addSub_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  addSub_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --addSub_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero971w972w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero973w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero973w974w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero971w & wire_altpriority_encoder20_w_lg_w_lg_zero973w974w);
	zero <= (wire_altpriority_encoder19_zero AND wire_altpriority_encoder20_zero);
	altpriority_encoder19 :  addSub_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder19_q,
		zero => wire_altpriority_encoder19_zero
	  );
	loop59 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero971w972w(i) <= wire_altpriority_encoder20_w_lg_zero971w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder20_w_lg_zero973w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop60;
	wire_altpriority_encoder20_w_lg_zero971w(0) <= NOT wire_altpriority_encoder20_zero;
	loop61 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero973w974w(i) <= wire_altpriority_encoder20_w_lg_zero973w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero971w972w(i);
	END GENERATE loop61;
	altpriority_encoder20 :  addSub_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --addSub_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero906w907w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero908w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero908w909w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder8_w_lg_zero906w & wire_altpriority_encoder8_w_lg_w_lg_zero908w909w);
	altpriority_encoder7 :  addSub_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder7_q
	  );
	loop62 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero906w907w(i) <= wire_altpriority_encoder8_w_lg_zero906w(0) AND wire_altpriority_encoder8_q(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder8_w_lg_zero908w(i) <= wire_altpriority_encoder8_zero AND wire_altpriority_encoder7_q(i);
	END GENERATE loop63;
	wire_altpriority_encoder8_w_lg_zero906w(0) <= NOT wire_altpriority_encoder8_zero;
	loop64 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero908w909w(i) <= wire_altpriority_encoder8_w_lg_zero908w(i) OR wire_altpriority_encoder8_w_lg_w_lg_zero906w907w(i);
	END GENERATE loop64;
	altpriority_encoder8 :  addSub_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder8_q,
		zero => wire_altpriority_encoder8_zero
	  );

 END RTL; --addSub_altpriority_encoder_qb6


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_nh8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_nh8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_nh8 IS

	 SIGNAL  wire_altpriority_encoder27_w_lg_w_data_range1018w1020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_w_data_range1018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altpriority_encoder27_w_lg_w_data_range1018w1020w(0) <= NOT wire_altpriority_encoder27_w_data_range1018w(0);
	q <= ( wire_altpriority_encoder27_w_lg_w_data_range1018w1020w);
	zero <= (NOT (data(0) OR data(1)));
	wire_altpriority_encoder27_w_data_range1018w(0) <= data(0);

 END RTL; --addSub_altpriority_encoder_nh8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_qh8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_qh8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_qh8 IS

	 SIGNAL  wire_altpriority_encoder27_w_lg_w_lg_zero1010w1011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_w_lg_zero1012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_w_lg_zero1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_w_lg_w_lg_zero1012w1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder27_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder28_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder28_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_nh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder27_zero & wire_altpriority_encoder27_w_lg_w_lg_zero1012w1013w);
	zero <= (wire_altpriority_encoder27_zero AND wire_altpriority_encoder28_zero);
	wire_altpriority_encoder27_w_lg_w_lg_zero1010w1011w(0) <= wire_altpriority_encoder27_w_lg_zero1010w(0) AND wire_altpriority_encoder27_q(0);
	wire_altpriority_encoder27_w_lg_zero1012w(0) <= wire_altpriority_encoder27_zero AND wire_altpriority_encoder28_q(0);
	wire_altpriority_encoder27_w_lg_zero1010w(0) <= NOT wire_altpriority_encoder27_zero;
	wire_altpriority_encoder27_w_lg_w_lg_zero1012w1013w(0) <= wire_altpriority_encoder27_w_lg_zero1012w(0) OR wire_altpriority_encoder27_w_lg_w_lg_zero1010w1011w(0);
	altpriority_encoder27 :  addSub_altpriority_encoder_nh8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder27_q,
		zero => wire_altpriority_encoder27_zero
	  );
	altpriority_encoder28 :  addSub_altpriority_encoder_nh8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder28_q,
		zero => wire_altpriority_encoder28_zero
	  );

 END RTL; --addSub_altpriority_encoder_qh8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_vh8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_vh8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_vh8 IS

	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1000w1001w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1002w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1002w1003w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder26_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder26_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_qh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder25_zero & wire_altpriority_encoder25_w_lg_w_lg_zero1002w1003w);
	zero <= (wire_altpriority_encoder25_zero AND wire_altpriority_encoder26_zero);
	loop65 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1000w1001w(i) <= wire_altpriority_encoder25_w_lg_zero1000w(0) AND wire_altpriority_encoder25_q(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder25_w_lg_zero1002w(i) <= wire_altpriority_encoder25_zero AND wire_altpriority_encoder26_q(i);
	END GENERATE loop66;
	wire_altpriority_encoder25_w_lg_zero1000w(0) <= NOT wire_altpriority_encoder25_zero;
	loop67 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1002w1003w(i) <= wire_altpriority_encoder25_w_lg_zero1002w(i) OR wire_altpriority_encoder25_w_lg_w_lg_zero1000w1001w(i);
	END GENERATE loop67;
	altpriority_encoder25 :  addSub_altpriority_encoder_qh8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder25_q,
		zero => wire_altpriority_encoder25_zero
	  );
	altpriority_encoder26 :  addSub_altpriority_encoder_qh8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder26_q,
		zero => wire_altpriority_encoder26_zero
	  );

 END RTL; --addSub_altpriority_encoder_vh8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_fj8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END addSub_altpriority_encoder_fj8;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_fj8 IS

	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero990w991w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero992w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero992w993w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder24_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder24_zero	:	STD_LOGIC;
	 COMPONENT  addSub_altpriority_encoder_vh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder23_zero & wire_altpriority_encoder23_w_lg_w_lg_zero992w993w);
	zero <= (wire_altpriority_encoder23_zero AND wire_altpriority_encoder24_zero);
	loop68 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero990w991w(i) <= wire_altpriority_encoder23_w_lg_zero990w(0) AND wire_altpriority_encoder23_q(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder23_w_lg_zero992w(i) <= wire_altpriority_encoder23_zero AND wire_altpriority_encoder24_q(i);
	END GENERATE loop69;
	wire_altpriority_encoder23_w_lg_zero990w(0) <= NOT wire_altpriority_encoder23_zero;
	loop70 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero992w993w(i) <= wire_altpriority_encoder23_w_lg_zero992w(i) OR wire_altpriority_encoder23_w_lg_w_lg_zero990w991w(i);
	END GENERATE loop70;
	altpriority_encoder23 :  addSub_altpriority_encoder_vh8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder23_q,
		zero => wire_altpriority_encoder23_zero
	  );
	altpriority_encoder24 :  addSub_altpriority_encoder_vh8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder24_q,
		zero => wire_altpriority_encoder24_zero
	  );

 END RTL; --addSub_altpriority_encoder_fj8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="YES" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_n28 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_n28;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_n28 IS

	 SIGNAL  wire_altpriority_encoder34_w_lg_w_data_range1052w1054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder34_w_data_range1052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altpriority_encoder34_w_lg_w_data_range1052w1054w(0) <= NOT wire_altpriority_encoder34_w_data_range1052w(0);
	q <= ( wire_altpriority_encoder34_w_lg_w_data_range1052w1054w);
	wire_altpriority_encoder34_w_data_range1052w(0) <= data(0);

 END RTL; --addSub_altpriority_encoder_n28

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_q28 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_q28;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_q28 IS

	 SIGNAL  wire_altpriority_encoder33_w_lg_w_lg_zero1045w1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder33_w_lg_zero1047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder33_w_lg_zero1045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder33_w_lg_w_lg_zero1047w1048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder33_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder33_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder34_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  addSub_altpriority_encoder_nh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_n28
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder33_zero & wire_altpriority_encoder33_w_lg_w_lg_zero1047w1048w);
	wire_altpriority_encoder33_w_lg_w_lg_zero1045w1046w(0) <= wire_altpriority_encoder33_w_lg_zero1045w(0) AND wire_altpriority_encoder33_q(0);
	wire_altpriority_encoder33_w_lg_zero1047w(0) <= wire_altpriority_encoder33_zero AND wire_altpriority_encoder34_q(0);
	wire_altpriority_encoder33_w_lg_zero1045w(0) <= NOT wire_altpriority_encoder33_zero;
	wire_altpriority_encoder33_w_lg_w_lg_zero1047w1048w(0) <= wire_altpriority_encoder33_w_lg_zero1047w(0) OR wire_altpriority_encoder33_w_lg_w_lg_zero1045w1046w(0);
	altpriority_encoder33 :  addSub_altpriority_encoder_nh8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder33_q,
		zero => wire_altpriority_encoder33_zero
	  );
	altpriority_encoder34 :  addSub_altpriority_encoder_n28
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder34_q
	  );

 END RTL; --addSub_altpriority_encoder_q28

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_v28 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_v28;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_v28 IS

	 SIGNAL  wire_altpriority_encoder31_w_lg_w_lg_zero1036w1037w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder31_w_lg_zero1038w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder31_w_lg_zero1036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder31_w_lg_w_lg_zero1038w1039w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder31_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder31_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder32_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 COMPONENT  addSub_altpriority_encoder_qh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_q28
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder31_zero & wire_altpriority_encoder31_w_lg_w_lg_zero1038w1039w);
	loop71 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder31_w_lg_w_lg_zero1036w1037w(i) <= wire_altpriority_encoder31_w_lg_zero1036w(0) AND wire_altpriority_encoder31_q(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder31_w_lg_zero1038w(i) <= wire_altpriority_encoder31_zero AND wire_altpriority_encoder32_q(i);
	END GENERATE loop72;
	wire_altpriority_encoder31_w_lg_zero1036w(0) <= NOT wire_altpriority_encoder31_zero;
	loop73 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder31_w_lg_w_lg_zero1038w1039w(i) <= wire_altpriority_encoder31_w_lg_zero1038w(i) OR wire_altpriority_encoder31_w_lg_w_lg_zero1036w1037w(i);
	END GENERATE loop73;
	altpriority_encoder31 :  addSub_altpriority_encoder_qh8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder31_q,
		zero => wire_altpriority_encoder31_zero
	  );
	altpriority_encoder32 :  addSub_altpriority_encoder_q28
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder32_q
	  );

 END RTL; --addSub_altpriority_encoder_v28

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_f48 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_f48;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_f48 IS

	 SIGNAL  wire_altpriority_encoder29_w_lg_w_lg_zero1027w1028w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder29_w_lg_zero1029w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder29_w_lg_zero1027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder29_w_lg_w_lg_zero1029w1030w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder29_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder29_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder30_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 COMPONENT  addSub_altpriority_encoder_vh8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_v28
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder29_zero & wire_altpriority_encoder29_w_lg_w_lg_zero1029w1030w);
	loop74 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder29_w_lg_w_lg_zero1027w1028w(i) <= wire_altpriority_encoder29_w_lg_zero1027w(0) AND wire_altpriority_encoder29_q(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder29_w_lg_zero1029w(i) <= wire_altpriority_encoder29_zero AND wire_altpriority_encoder30_q(i);
	END GENERATE loop75;
	wire_altpriority_encoder29_w_lg_zero1027w(0) <= NOT wire_altpriority_encoder29_zero;
	loop76 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder29_w_lg_w_lg_zero1029w1030w(i) <= wire_altpriority_encoder29_w_lg_zero1029w(i) OR wire_altpriority_encoder29_w_lg_w_lg_zero1027w1028w(i);
	END GENERATE loop76;
	altpriority_encoder29 :  addSub_altpriority_encoder_vh8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder29_q,
		zero => wire_altpriority_encoder29_zero
	  );
	altpriority_encoder30 :  addSub_altpriority_encoder_v28
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder30_q
	  );

 END RTL; --addSub_altpriority_encoder_f48

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altpriority_encoder_e48 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END addSub_altpriority_encoder_e48;

 ARCHITECTURE RTL OF addSub_altpriority_encoder_e48 IS

	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero981w982w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero983w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero983w984w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  addSub_altpriority_encoder_fj8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_f48
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder21_zero & wire_altpriority_encoder21_w_lg_w_lg_zero983w984w);
	loop77 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero981w982w(i) <= wire_altpriority_encoder21_w_lg_zero981w(0) AND wire_altpriority_encoder21_q(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder21_w_lg_zero983w(i) <= wire_altpriority_encoder21_zero AND wire_altpriority_encoder22_q(i);
	END GENERATE loop78;
	wire_altpriority_encoder21_w_lg_zero981w(0) <= NOT wire_altpriority_encoder21_zero;
	loop79 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero983w984w(i) <= wire_altpriority_encoder21_w_lg_zero983w(i) OR wire_altpriority_encoder21_w_lg_w_lg_zero981w982w(i);
	END GENERATE loop79;
	altpriority_encoder21 :  addSub_altpriority_encoder_fj8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );
	altpriority_encoder22 :  addSub_altpriority_encoder_f48
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder22_q
	  );

 END RTL; --addSub_altpriority_encoder_e48

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 14 lpm_compare 1 reg 283 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  addSub_altfp_add_sub_kdk IS 
	 PORT 
	 ( 
		 add_sub	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END addSub_altfp_add_sub_kdk;

 ARCHITECTURE RTL OF addSub_altfp_add_sub_kdk IS

	 SIGNAL  wire_lbarrel_shift_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_data	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_rbarrel_shift_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_leading_zeroes_cnt_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_leading_zeroes_cnt_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_trailing_zeros_cnt_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_trailing_zeros_cnt_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 add_sub_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 both_inputs_are_infinite_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 data_exp_dffe1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dataa_man_dffe1	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dataa_sign_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_man_dffe1	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_sign_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 denormal_res_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 denormal_res_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_adj_dffe21	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_out_dffe5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_res_dffe2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_res_dffe21	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_res_dffe3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_res_dffe4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_output_sign_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_res_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_res_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_magnitude_sub_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_magnitude_sub_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_magnitude_sub_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_magnitude_sub_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_magnitude_sub_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinite_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_add_sub_res_mag_dffe21	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_add_sub_res_sign_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe31	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_leading_zeros_dffe31	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_out_dffe5	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_res_dffe4	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_res_is_not_zero_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_res_is_not_zero_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_res_is_not_zero_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 need_complement_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_bit_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_bit_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 round_bit_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rounded_res_infinity_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_out_dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_res_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_res_dffe4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_bit_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_bit_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_bit_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_bit_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_bit_dffe31	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_man_sign_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_man_sign_dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_man_2comp_res_lower_w_lg_w_lg_cout381w382w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_2comp_res_lower_w_lg_cout380w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_2comp_res_lower_w_lg_cout381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_2comp_res_lower_w_lg_w_lg_w_lg_cout381w382w383w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_2comp_res_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_man_2comp_res_lower_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_man_2comp_res_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_man_2comp_res_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_lower_w_lg_w_lg_cout368w369w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_lower_w_lg_cout367w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_lower_w_lg_cout368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_lower_w_lg_w_lg_w_lg_cout368w369w370w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_man_add_sub_lower_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_add_sub_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_lower_w_lg_w_lg_cout594w595w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_lower_w_lg_cout593w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_lower_w_lg_cout594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_lower_w_lg_w_lg_w_lg_cout594w595w596w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_man_res_rounding_add_sub_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_man_res_rounding_add_sub_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_trailing_zeros_limit_comparator_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_dataa_sign_dffe1_wo345w349w350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w411w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_sign_dffe1_wo342w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_force_zero_w648w649w650w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_force_zero_w648w649w659w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_sign_dffe1_wo345w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_sign_dffe1_wo345w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_denormal_result_w572w573w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w324w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w331w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w317w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_amb_mux_w275w278w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_amb_mux_w275w276w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_infinity_w643w653w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_infinity_w643w662w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_infinity_w643w668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_nan_w644w656w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_nan_w644w665w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w243w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w234w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_dataa_infinite_dffe11_wo246w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w262w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w253w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_datab_infinite_dffe11_wo265w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_datab_infinite_dffe15_wo339w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_res_not_zero_dffe26_wo517w518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w292w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w397w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w426w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_man_add_sub_w_range386w389w392w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_w601w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_zero_w648w651w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_zero_w648w660w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_dataa_sign_dffe1_wo351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dataa_sign_dffe1_wo342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_dffe15_wo330w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_dffe15_wo323w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_dffe15_wo314w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_w279w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_w273w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_infinity_w654w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_infinity_w663w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_nan_w657w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_nan_w666w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_infinite_dffe15_wo338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_need_complement_dffe22_wo390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range17w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range27w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range37w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range47w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range57w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range67w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range77w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range20w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range30w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range40w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range50w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range60w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range70w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range80w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_all_one_w_range84w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_all_one_w_range86w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w293w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range554w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range557w558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range559w560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range563w564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range565w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range567w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_max_w_range569w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range615w618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range619w621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range622w624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range625w627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range628w630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range631w633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_rounded_res_max_w_range634w636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w398w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w428w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_w_range386w393w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_rounding_add_sub_w_range599w603w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_zero_w648w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_aligned_datab_sign_dffe15_wo336w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_sub_dffe1_wo344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_sub_dffe25_wo505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_sub_w2356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dataa_sign_dffe1_wo345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_datab_sign_dffe1_wo348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_result_w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_dffe15_wo316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_amb_mux_w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_infinity_w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_nan_w644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_zero_w642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_dataa_denormal_dffe11_wo233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_dataa_infinite_dffe11_wo246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_dataa_zero_dffe11_wo245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_denormal_dffe11_wo252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_infinite_dffe11_wo265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_infinite_dffe15_wo339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_zero_dffe11_wo264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_res_is_not_zero_dffe4_wo641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_res_not_zero_dffe26_wo517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_need_complement_dffe22_wo387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sticky_bit_dffe1_wo357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_adjustment2_add_sub_w_range525w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_not_zero_w_range215w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range401w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_add_sub_w_range386w389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_not_zero_w_range218w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_rounding_add_sub_w_range599w600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_force_zero_w648w651w652w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_force_zero_w648w660w661w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_infinity_w654w655w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_force_infinity_w663w664w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_force_zero_w648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sticky_bit_dffe27_wo416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range147w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range153w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range183w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range189w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range195w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range87w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range17w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range27w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range37w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range47w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range77w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range156w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range162w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range174w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range198w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range20w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range30w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range40w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range80w81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_diff_abs_exceed_max_w_range282w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_diff_abs_exceed_max_w_range286w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range530w533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range534w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range537w539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range540w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range543w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range546w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range549w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_not_zero_w_range552w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range431w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range462w464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range465w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range468w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range471w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range474w476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range477w479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range480w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range483w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range486w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range489w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range435w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range492w494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range495w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range498w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range501w503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range438w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range441w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range444w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range447w449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range450w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range453w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range456w458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_not_zero_w2_range459w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_aligned_datab_sign_dffe15_wo336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_sub_dffe11_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe11_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe12_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe12_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe13_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe13_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe14_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe14_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe15_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe15_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe1_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe1_wo :	STD_LOGIC;
	 SIGNAL  add_sub_dffe25_wi :	STD_LOGIC;
	 SIGNAL  add_sub_dffe25_wo :	STD_LOGIC;
	 SIGNAL  add_sub_w2 :	STD_LOGIC;
	 SIGNAL  adder_upper_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe12_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe12_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe13_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe13_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe14_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe14_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe15_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_dffe15_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_exp_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe12_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe12_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe13_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe13_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe14_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe14_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe15_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe15_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_dffe15_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_dataa_man_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  aligned_dataa_sign_dffe12_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe12_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe13_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe13_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe14_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe14_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe15_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe15_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_w :	STD_LOGIC;
	 SIGNAL  aligned_datab_exp_dffe12_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe12_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe13_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe13_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe14_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe14_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe15_wi :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_dffe15_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_exp_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe12_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe12_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe13_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe13_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe14_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe14_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe15_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe15_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_dffe15_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  aligned_datab_man_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  aligned_datab_sign_dffe12_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe12_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe13_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe13_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe14_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe14_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe15_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe15_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_w :	STD_LOGIC;
	 SIGNAL  borrow_w :	STD_LOGIC;
	 SIGNAL  both_inputs_are_infinite_dffe1_wi :	STD_LOGIC;
	 SIGNAL  both_inputs_are_infinite_dffe1_wo :	STD_LOGIC;
	 SIGNAL  both_inputs_are_infinite_dffe25_wi :	STD_LOGIC;
	 SIGNAL  both_inputs_are_infinite_dffe25_wo :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  data_exp_dffe1_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  data_exp_dffe1_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  dataa_dffe11_wi :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dataa_dffe11_wo :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dataa_man_dffe1_wi :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  dataa_man_dffe1_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  dataa_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  dataa_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  dataa_sign_dffe25_wi :	STD_LOGIC;
	 SIGNAL  dataa_sign_dffe25_wo :	STD_LOGIC;
	 SIGNAL  datab_dffe11_wi :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  datab_dffe11_wo :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  datab_man_dffe1_wi :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  datab_man_dffe1_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  datab_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  datab_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  denormal_flag_w :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe32_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe32_wo :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe33_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe33_wo :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe3_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe3_wo :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe41_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe41_wo :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe42_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe42_wo :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe4_wi :	STD_LOGIC;
	 SIGNAL  denormal_res_dffe4_wo :	STD_LOGIC;
	 SIGNAL  denormal_result_w :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_adj_0pads :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  exp_adj_dffe21_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adj_dffe21_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adj_dffe23_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adj_dffe23_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adj_dffe26_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adj_dffe26_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adjust_by_add1 :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adjust_by_add2 :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_adjustment2_add_sub_dataa_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_adjustment2_add_sub_datab_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_adjustment2_add_sub_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_adjustment_add_sub_dataa_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_adjustment_add_sub_datab_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_adjustment_add_sub_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_all_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_all_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_amb_mux_dffe13_wi :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_dffe13_wo :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_dffe14_wi :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_dffe14_wo :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_dffe15_wi :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_dffe15_wo :	STD_LOGIC;
	 SIGNAL  exp_amb_mux_w :	STD_LOGIC;
	 SIGNAL  exp_amb_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_b_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_bma_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_diff_abs_exceed_max_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  exp_diff_abs_max_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  exp_diff_abs_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_intermediate_res_dffe41_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_intermediate_res_dffe41_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_intermediate_res_dffe42_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_intermediate_res_dffe42_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_intermediate_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_out_dffe5_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_out_dffe5_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe21_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe21_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe22_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe22_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe23_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe23_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe25_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe25_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe26_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe26_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe27_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe27_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe2_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe2_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe32_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe32_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe33_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe33_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe3_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe3_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe4_wi :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_dffe4_wo :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_max_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_not_zero_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_res_rounding_adder_dataa_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_res_rounding_adder_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_rounded_res_infinity_w :	STD_LOGIC;
	 SIGNAL  exp_rounded_res_max_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_rounded_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_rounding_adjustment_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_value :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  force_infinity_w :	STD_LOGIC;
	 SIGNAL  force_nan_w :	STD_LOGIC;
	 SIGNAL  force_zero_w :	STD_LOGIC;
	 SIGNAL  guard_bit_dffe3_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe21_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe21_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe22_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe22_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe23_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe23_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe25_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe25_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe26_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe26_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe27_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe27_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe2_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe2_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe31_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe31_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe32_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe32_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe33_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe33_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe3_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe3_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe41_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe41_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe42_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe42_wo :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe4_wi :	STD_LOGIC;
	 SIGNAL  infinite_output_sign_dffe4_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dff32_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dff32_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dff33_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dff33_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe3_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe3_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe41_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe41_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe42_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe42_wo :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe4_wi :	STD_LOGIC;
	 SIGNAL  infinite_res_dffe4_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe21_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe21_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe22_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe22_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe23_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe23_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe26_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe26_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe27_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe27_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe2_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe2_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe31_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe31_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe32_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe32_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe33_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe33_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe3_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe3_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe41_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe41_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe42_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe42_wo :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe4_wi :	STD_LOGIC;
	 SIGNAL  infinity_magnitude_sub_dffe4_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_denormal_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_denormal_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_denormal_w :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe12_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe12_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe13_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe13_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe14_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe14_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe15_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_dffe15_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_infinite_w :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe12_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe12_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_w :	STD_LOGIC;
	 SIGNAL  input_dataa_zero_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_zero_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_zero_w :	STD_LOGIC;
	 SIGNAL  input_datab_denormal_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_datab_denormal_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_datab_denormal_w :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe12_wi :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe12_wo :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe13_wi :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe13_wo :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe14_wi :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe14_wo :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe15_wi :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_dffe15_wo :	STD_LOGIC;
	 SIGNAL  input_datab_infinite_w :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe12_wi :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe12_wo :	STD_LOGIC;
	 SIGNAL  input_datab_nan_w :	STD_LOGIC;
	 SIGNAL  input_datab_zero_dffe11_wi :	STD_LOGIC;
	 SIGNAL  input_datab_zero_dffe11_wo :	STD_LOGIC;
	 SIGNAL  input_datab_zero_w :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe1_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe1_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe21_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe21_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe22_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe22_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe23_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe23_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe25_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe25_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe26_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe26_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe27_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe27_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe31_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe31_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe32_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe32_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe33_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe33_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe3_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe3_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe41_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe41_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe42_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe42_wo :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe4_wi :	STD_LOGIC;
	 SIGNAL  input_is_infinite_dffe4_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe13_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe13_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe14_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe14_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe15_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe15_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe1_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe1_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe21_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe21_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe22_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe22_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe23_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe23_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe25_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe25_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe26_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe26_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe27_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe27_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe31_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe31_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe32_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe32_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe33_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe33_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe3_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe3_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe41_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe41_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe42_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe42_wo :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe4_wi :	STD_LOGIC;
	 SIGNAL  input_is_nan_dffe4_wo :	STD_LOGIC;
	 SIGNAL  man_2comp_res_dataa_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_2comp_res_datab_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_2comp_res_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_a_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_add_sub_dataa_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_add_sub_datab_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe21_wi :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe21_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe23_wi :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe23_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe26_wi :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe26_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe27_wi :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_dffe27_wo :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_add_sub_res_mag_w2 :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_add_sub_res_sign_dffe21_wo :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe23_wi :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe23_wo :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe26_wi :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe26_wo :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe27_wi :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_dffe27_wo :	STD_LOGIC;
	 SIGNAL  man_add_sub_res_sign_w2 :	STD_LOGIC;
	 SIGNAL  man_add_sub_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  man_all_zeros_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_dffe31_wo :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_intermediate_res_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_leading_zeros_cnt_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  man_leading_zeros_dffe31_wi :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  man_leading_zeros_dffe31_wo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  man_nan_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_out_dffe5_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_out_dffe5_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_dffe4_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_dffe4_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_is_not_zero_dffe31_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe31_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe32_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe32_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe33_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe33_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe3_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe3_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe41_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe41_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe42_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe42_wo :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe4_wi :	STD_LOGIC;
	 SIGNAL  man_res_is_not_zero_dffe4_wo :	STD_LOGIC;
	 SIGNAL  man_res_mag_w2 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_res_not_zero_dffe23_wi :	STD_LOGIC;
	 SIGNAL  man_res_not_zero_dffe23_wo :	STD_LOGIC;
	 SIGNAL  man_res_not_zero_dffe26_wi :	STD_LOGIC;
	 SIGNAL  man_res_not_zero_dffe26_wo :	STD_LOGIC;
	 SIGNAL  man_res_not_zero_w2 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_res_rounding_add_sub_datab_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_res_rounding_add_sub_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  man_res_w3 :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_rounded_res_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_rounding_add_value_w :	STD_LOGIC;
	 SIGNAL  man_smaller_dffe13_wi :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_smaller_dffe13_wo :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_smaller_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  need_complement_dffe22_wi :	STD_LOGIC;
	 SIGNAL  need_complement_dffe22_wo :	STD_LOGIC;
	 SIGNAL  need_complement_dffe2_wi :	STD_LOGIC;
	 SIGNAL  need_complement_dffe2_wo :	STD_LOGIC;
	 SIGNAL  pos_sign_bit_ext :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  priority_encoder_1pads_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  round_bit_dffe21_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe21_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe23_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe23_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe26_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe26_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe31_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe31_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe32_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe32_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe33_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe33_wo :	STD_LOGIC;
	 SIGNAL  round_bit_dffe3_wi :	STD_LOGIC;
	 SIGNAL  round_bit_dffe3_wo :	STD_LOGIC;
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  rounded_res_infinity_dffe4_wi :	STD_LOGIC;
	 SIGNAL  rounded_res_infinity_dffe4_wo :	STD_LOGIC;
	 SIGNAL  rshift_distance_dffe13_wi :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_dffe13_wo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_dffe14_wi :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_dffe14_wo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_dffe15_wi :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_dffe15_wo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rshift_distance_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  sign_dffe31_wi :	STD_LOGIC;
	 SIGNAL  sign_dffe31_wo :	STD_LOGIC;
	 SIGNAL  sign_dffe32_wi :	STD_LOGIC;
	 SIGNAL  sign_dffe32_wo :	STD_LOGIC;
	 SIGNAL  sign_dffe33_wi :	STD_LOGIC;
	 SIGNAL  sign_dffe33_wo :	STD_LOGIC;
	 SIGNAL  sign_out_dffe5_wi :	STD_LOGIC;
	 SIGNAL  sign_out_dffe5_wo :	STD_LOGIC;
	 SIGNAL  sign_res_dffe3_wi :	STD_LOGIC;
	 SIGNAL  sign_res_dffe3_wo :	STD_LOGIC;
	 SIGNAL  sign_res_dffe41_wi :	STD_LOGIC;
	 SIGNAL  sign_res_dffe41_wo :	STD_LOGIC;
	 SIGNAL  sign_res_dffe42_wi :	STD_LOGIC;
	 SIGNAL  sign_res_dffe42_wo :	STD_LOGIC;
	 SIGNAL  sign_res_dffe4_wi :	STD_LOGIC;
	 SIGNAL  sign_res_dffe4_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_cnt_dataa_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_cnt_datab_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_cnt_res_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_dffe1_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe1_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe21_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe21_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe22_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe22_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe23_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe23_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe25_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe25_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe26_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe26_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe27_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe27_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe2_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe2_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe31_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe31_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe32_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe32_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe33_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe33_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe3_wi :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe3_wo :	STD_LOGIC;
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  trailing_zeros_limit_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  zero_man_sign_dffe21_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe21_wo :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe22_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe22_wo :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe23_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe23_wo :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe26_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe26_wo :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe27_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe27_wo :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe2_wi :	STD_LOGIC;
	 SIGNAL  zero_man_sign_dffe2_wo :	STD_LOGIC;
	 SIGNAL  wire_w_aligned_dataa_exp_dffe15_wo_range315w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_aligned_datab_exp_dffe15_wo_range313w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_dffe11_wo_range242w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_dataa_dffe11_wo_range232w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_dffe11_wo_range261w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_datab_dffe11_wo_range251w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range571w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_adjustment2_add_sub_w_range525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_amb_w_range274w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bma_w_range272w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_exceed_max_w_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_exceed_max_w_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_exceed_max_w_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_w_range290w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_w_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_diff_abs_w_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_max_w_range569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_not_zero_w_range552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_max_w_range634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_rounded_res_w_range635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe21_wo_range454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe27_wo_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe27_wo_range425w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe27_wo_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe27_wo_range427w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_res_mag_dffe27_wo_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_add_sub_w_range386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_not_zero_w2_range459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_rounding_add_sub_w_range598w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_man_res_rounding_add_sub_w_range602w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_man_res_rounding_add_sub_w_range599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  addSub_altbarrel_shift_35e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altbarrel_shift_olb
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  addSub_altpriority_encoder_e48
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_w_lg_w_lg_w_lg_dataa_sign_dffe1_wo345w349w350w(0) <= wire_w_lg_w_lg_dataa_sign_dffe1_wo345w349w(0) AND add_sub_dffe1_wo;
	wire_w248w(0) <= wire_w_lg_w_lg_input_dataa_infinite_dffe11_wo246w247w(0) AND wire_w_lg_input_dataa_zero_dffe11_wo245w(0);
	wire_w267w(0) <= wire_w_lg_w_lg_input_datab_infinite_dffe11_wo265w266w(0) AND wire_w_lg_input_datab_zero_dffe11_wo264w(0);
	wire_w_lg_w411w421w(0) <= wire_w411w(0) AND sticky_bit_dffe27_wo;
	wire_w_lg_w_lg_dataa_sign_dffe1_wo342w343w(0) <= wire_w_lg_dataa_sign_dffe1_wo342w(0) AND add_sub_dffe1_wo;
	loop80 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_force_zero_w648w649w650w(i) <= wire_w_lg_w_lg_force_zero_w648w649w(0) AND exp_res_dffe4_wo(i);
	END GENERATE loop80;
	loop81 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_force_zero_w648w649w659w(i) <= wire_w_lg_w_lg_force_zero_w648w649w(0) AND man_res_dffe4_wo(i);
	END GENERATE loop81;
	wire_w_lg_w_lg_dataa_sign_dffe1_wo345w349w(0) <= wire_w_lg_dataa_sign_dffe1_wo345w(0) AND wire_w_lg_datab_sign_dffe1_wo348w(0);
	wire_w_lg_w_lg_dataa_sign_dffe1_wo345w346w(0) <= wire_w_lg_dataa_sign_dffe1_wo345w(0) AND datab_sign_dffe1_wo;
	loop82 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_denormal_result_w572w573w(i) <= wire_w_lg_denormal_result_w572w(0) AND wire_w_exp_adjustment2_add_sub_w_range571w(i);
	END GENERATE loop82;
	loop83 : FOR i IN 0 TO 25 GENERATE 
		wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w324w(i) <= wire_w_lg_exp_amb_mux_dffe15_wo316w(0) AND aligned_dataa_man_dffe15_w(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 25 GENERATE 
		wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w331w(i) <= wire_w_lg_exp_amb_mux_dffe15_wo316w(0) AND wire_rbarrel_shift_result(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w317w(i) <= wire_w_lg_exp_amb_mux_dffe15_wo316w(0) AND wire_w_aligned_dataa_exp_dffe15_wo_range315w(i);
	END GENERATE loop85;
	loop86 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_w_lg_exp_amb_mux_w275w278w(i) <= wire_w_lg_exp_amb_mux_w275w(0) AND aligned_datab_man_dffe12_wo(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_exp_amb_mux_w275w276w(i) <= wire_w_lg_exp_amb_mux_w275w(0) AND wire_w_exp_amb_w_range274w(i);
	END GENERATE loop87;
	loop88 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_force_infinity_w643w653w(i) <= wire_w_lg_force_infinity_w643w(0) AND wire_w_lg_w_lg_w_lg_force_zero_w648w651w652w(i);
	END GENERATE loop88;
	loop89 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_force_infinity_w643w662w(i) <= wire_w_lg_force_infinity_w643w(0) AND wire_w_lg_w_lg_w_lg_force_zero_w648w660w661w(i);
	END GENERATE loop89;
	wire_w_lg_w_lg_force_infinity_w643w668w(0) <= wire_w_lg_force_infinity_w643w(0) AND sign_res_dffe4_wo;
	loop90 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_force_nan_w644w656w(i) <= wire_w_lg_force_nan_w644w(0) AND wire_w_lg_w_lg_force_infinity_w654w655w(i);
	END GENERATE loop90;
	loop91 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_force_nan_w644w665w(i) <= wire_w_lg_force_nan_w644w(0) AND wire_w_lg_w_lg_force_infinity_w663w664w(i);
	END GENERATE loop91;
	loop92 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w243w(i) <= wire_w_lg_input_dataa_denormal_dffe11_wo233w(0) AND wire_w_dataa_dffe11_wo_range242w(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w234w(i) <= wire_w_lg_input_dataa_denormal_dffe11_wo233w(0) AND wire_w_dataa_dffe11_wo_range232w(i);
	END GENERATE loop93;
	wire_w_lg_w_lg_input_dataa_infinite_dffe11_wo246w247w(0) <= wire_w_lg_input_dataa_infinite_dffe11_wo246w(0) AND wire_w_lg_input_dataa_denormal_dffe11_wo233w(0);
	loop94 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w262w(i) <= wire_w_lg_input_datab_denormal_dffe11_wo252w(0) AND wire_w_datab_dffe11_wo_range261w(i);
	END GENERATE loop94;
	loop95 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w253w(i) <= wire_w_lg_input_datab_denormal_dffe11_wo252w(0) AND wire_w_datab_dffe11_wo_range251w(i);
	END GENERATE loop95;
	wire_w_lg_w_lg_input_datab_infinite_dffe11_wo265w266w(0) <= wire_w_lg_input_datab_infinite_dffe11_wo265w(0) AND wire_w_lg_input_datab_denormal_dffe11_wo252w(0);
	wire_w_lg_w_lg_input_datab_infinite_dffe15_wo339w340w(0) <= wire_w_lg_input_datab_infinite_dffe15_wo339w(0) AND aligned_dataa_sign_dffe15_wo;
	wire_w_lg_w_lg_man_res_not_zero_dffe26_wo517w518w(0) <= wire_w_lg_man_res_not_zero_dffe26_wo517w(0) AND zero_man_sign_dffe26_wo;
	loop96 : FOR i IN 0 TO 4 GENERATE 
		wire_w292w(i) <= wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w291w(0) AND wire_w_exp_diff_abs_w_range290w(i);
	END GENERATE loop96;
	wire_w411w(0) <= wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) AND wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range401w404w(0);
	loop97 : FOR i IN 0 TO 1 GENERATE 
		wire_w397w(i) <= wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) AND exp_adjust_by_add1(i);
	END GENERATE loop97;
	loop98 : FOR i IN 0 TO 25 GENERATE 
		wire_w426w(i) <= wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) AND wire_w_man_add_sub_res_mag_dffe27_wo_range425w(i);
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 27 GENERATE 
		wire_w_lg_w_lg_w_man_add_sub_w_range386w389w392w(i) <= wire_w_lg_w_man_add_sub_w_range386w389w(0) AND man_add_sub_w(i);
	END GENERATE loop99;
	loop100 : FOR i IN 0 TO 22 GENERATE 
		wire_w601w(i) <= wire_w_lg_w_man_res_rounding_add_sub_w_range599w600w(0) AND wire_w_man_res_rounding_add_sub_w_range598w(i);
	END GENERATE loop100;
	loop101 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_force_zero_w648w651w(i) <= wire_w_lg_force_zero_w648w(0) AND exp_all_zeros_w(i);
	END GENERATE loop101;
	loop102 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_force_zero_w648w660w(i) <= wire_w_lg_force_zero_w648w(0) AND man_all_zeros_w(i);
	END GENERATE loop102;
	wire_w_lg_dataa_sign_dffe1_wo351w(0) <= dataa_sign_dffe1_wo AND wire_w_lg_datab_sign_dffe1_wo348w(0);
	wire_w_lg_dataa_sign_dffe1_wo342w(0) <= dataa_sign_dffe1_wo AND datab_sign_dffe1_wo;
	loop103 : FOR i IN 0 TO 25 GENERATE 
		wire_w_lg_exp_amb_mux_dffe15_wo330w(i) <= exp_amb_mux_dffe15_wo AND aligned_datab_man_dffe15_w(i);
	END GENERATE loop103;
	loop104 : FOR i IN 0 TO 25 GENERATE 
		wire_w_lg_exp_amb_mux_dffe15_wo323w(i) <= exp_amb_mux_dffe15_wo AND wire_rbarrel_shift_result(i);
	END GENERATE loop104;
	loop105 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_exp_amb_mux_dffe15_wo314w(i) <= exp_amb_mux_dffe15_wo AND wire_w_aligned_datab_exp_dffe15_wo_range313w(i);
	END GENERATE loop105;
	loop106 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_exp_amb_mux_w279w(i) <= exp_amb_mux_w AND aligned_dataa_man_dffe12_wo(i);
	END GENERATE loop106;
	loop107 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_exp_amb_mux_w273w(i) <= exp_amb_mux_w AND wire_w_exp_bma_w_range272w(i);
	END GENERATE loop107;
	loop108 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_force_infinity_w654w(i) <= force_infinity_w AND exp_all_ones_w(i);
	END GENERATE loop108;
	loop109 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_force_infinity_w663w(i) <= force_infinity_w AND man_all_zeros_w(i);
	END GENERATE loop109;
	loop110 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_force_nan_w657w(i) <= force_nan_w AND exp_all_ones_w(i);
	END GENERATE loop110;
	loop111 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_force_nan_w666w(i) <= force_nan_w AND man_nan_w(i);
	END GENERATE loop111;
	wire_w_lg_input_datab_infinite_dffe15_wo338w(0) <= input_datab_infinite_dffe15_wo AND wire_w_lg_w_lg_aligned_datab_sign_dffe15_wo336w337w(0);
	wire_w_lg_need_complement_dffe22_wo390w(0) <= need_complement_dffe22_wo AND wire_w_lg_w_man_add_sub_w_range386w389w(0);
	wire_w_lg_w_dataa_range17w23w(0) <= wire_w_dataa_range17w(0) AND wire_w_exp_a_all_one_w_range7w(0);
	wire_w_lg_w_dataa_range27w33w(0) <= wire_w_dataa_range27w(0) AND wire_w_exp_a_all_one_w_range24w(0);
	wire_w_lg_w_dataa_range37w43w(0) <= wire_w_dataa_range37w(0) AND wire_w_exp_a_all_one_w_range34w(0);
	wire_w_lg_w_dataa_range47w53w(0) <= wire_w_dataa_range47w(0) AND wire_w_exp_a_all_one_w_range44w(0);
	wire_w_lg_w_dataa_range57w63w(0) <= wire_w_dataa_range57w(0) AND wire_w_exp_a_all_one_w_range54w(0);
	wire_w_lg_w_dataa_range67w73w(0) <= wire_w_dataa_range67w(0) AND wire_w_exp_a_all_one_w_range64w(0);
	wire_w_lg_w_dataa_range77w83w(0) <= wire_w_dataa_range77w(0) AND wire_w_exp_a_all_one_w_range74w(0);
	wire_w_lg_w_datab_range20w25w(0) <= wire_w_datab_range20w(0) AND wire_w_exp_b_all_one_w_range9w(0);
	wire_w_lg_w_datab_range30w35w(0) <= wire_w_datab_range30w(0) AND wire_w_exp_b_all_one_w_range26w(0);
	wire_w_lg_w_datab_range40w45w(0) <= wire_w_datab_range40w(0) AND wire_w_exp_b_all_one_w_range36w(0);
	wire_w_lg_w_datab_range50w55w(0) <= wire_w_datab_range50w(0) AND wire_w_exp_b_all_one_w_range46w(0);
	wire_w_lg_w_datab_range60w65w(0) <= wire_w_datab_range60w(0) AND wire_w_exp_b_all_one_w_range56w(0);
	wire_w_lg_w_datab_range70w75w(0) <= wire_w_datab_range70w(0) AND wire_w_exp_b_all_one_w_range66w(0);
	wire_w_lg_w_datab_range80w85w(0) <= wire_w_datab_range80w(0) AND wire_w_exp_b_all_one_w_range76w(0);
	wire_w_lg_w_exp_a_all_one_w_range84w220w(0) <= wire_w_exp_a_all_one_w_range84w(0) AND wire_w_lg_w_man_a_not_zero_w_range215w219w(0);
	wire_w_lg_w_exp_b_all_one_w_range86w226w(0) <= wire_w_exp_b_all_one_w_range86w(0) AND wire_w_lg_w_man_b_not_zero_w_range218w225w(0);
	loop112 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w293w(i) <= wire_w_exp_diff_abs_exceed_max_w_range289w(0) AND exp_diff_abs_max_w(i);
	END GENERATE loop112;
	wire_w_lg_w_exp_res_max_w_range554w556w(0) <= wire_w_exp_res_max_w_range554w(0) AND wire_w_exp_adjustment2_add_sub_w_range532w(0);
	wire_w_lg_w_exp_res_max_w_range557w558w(0) <= wire_w_exp_res_max_w_range557w(0) AND wire_w_exp_adjustment2_add_sub_w_range535w(0);
	wire_w_lg_w_exp_res_max_w_range559w560w(0) <= wire_w_exp_res_max_w_range559w(0) AND wire_w_exp_adjustment2_add_sub_w_range538w(0);
	wire_w_lg_w_exp_res_max_w_range561w562w(0) <= wire_w_exp_res_max_w_range561w(0) AND wire_w_exp_adjustment2_add_sub_w_range541w(0);
	wire_w_lg_w_exp_res_max_w_range563w564w(0) <= wire_w_exp_res_max_w_range563w(0) AND wire_w_exp_adjustment2_add_sub_w_range544w(0);
	wire_w_lg_w_exp_res_max_w_range565w566w(0) <= wire_w_exp_res_max_w_range565w(0) AND wire_w_exp_adjustment2_add_sub_w_range547w(0);
	wire_w_lg_w_exp_res_max_w_range567w568w(0) <= wire_w_exp_res_max_w_range567w(0) AND wire_w_exp_adjustment2_add_sub_w_range550w(0);
	wire_w_lg_w_exp_res_max_w_range569w575w(0) <= wire_w_exp_res_max_w_range569w(0) AND wire_w_lg_w_exp_adjustment2_add_sub_w_range525w574w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range615w618w(0) <= wire_w_exp_rounded_res_max_w_range615w(0) AND wire_w_exp_rounded_res_w_range617w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range619w621w(0) <= wire_w_exp_rounded_res_max_w_range619w(0) AND wire_w_exp_rounded_res_w_range620w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range622w624w(0) <= wire_w_exp_rounded_res_max_w_range622w(0) AND wire_w_exp_rounded_res_w_range623w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range625w627w(0) <= wire_w_exp_rounded_res_max_w_range625w(0) AND wire_w_exp_rounded_res_w_range626w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range628w630w(0) <= wire_w_exp_rounded_res_max_w_range628w(0) AND wire_w_exp_rounded_res_w_range629w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range631w633w(0) <= wire_w_exp_rounded_res_max_w_range631w(0) AND wire_w_exp_rounded_res_w_range632w(0);
	wire_w_lg_w_exp_rounded_res_max_w_range634w636w(0) <= wire_w_exp_rounded_res_max_w_range634w(0) AND wire_w_exp_rounded_res_w_range635w(0);
	wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w405w(0) <= wire_w_man_add_sub_res_mag_dffe27_wo_range395w(0) AND wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range401w404w(0);
	loop113 : FOR i IN 0 TO 1 GENERATE 
		wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w398w(i) <= wire_w_man_add_sub_res_mag_dffe27_wo_range395w(0) AND exp_adjust_by_add2(i);
	END GENERATE loop113;
	loop114 : FOR i IN 0 TO 25 GENERATE 
		wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w428w(i) <= wire_w_man_add_sub_res_mag_dffe27_wo_range395w(0) AND wire_w_man_add_sub_res_mag_dffe27_wo_range427w(i);
	END GENERATE loop114;
	loop115 : FOR i IN 0 TO 27 GENERATE 
		wire_w_lg_w_man_add_sub_w_range386w393w(i) <= wire_w_man_add_sub_w_range386w(0) AND man_2comp_res_w(i);
	END GENERATE loop115;
	loop116 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_man_res_rounding_add_sub_w_range599w603w(i) <= wire_w_man_res_rounding_add_sub_w_range599w(0) AND wire_w_man_res_rounding_add_sub_w_range602w(i);
	END GENERATE loop116;
	wire_w_lg_w_lg_force_zero_w648w649w(0) <= NOT wire_w_lg_force_zero_w648w(0);
	wire_w_lg_w_lg_aligned_datab_sign_dffe15_wo336w337w(0) <= NOT wire_w_lg_aligned_datab_sign_dffe15_wo336w(0);
	wire_w_lg_add_sub_dffe1_wo344w(0) <= NOT add_sub_dffe1_wo;
	wire_w_lg_add_sub_dffe25_wo505w(0) <= NOT add_sub_dffe25_wo;
	wire_w_lg_add_sub_w2356w(0) <= NOT add_sub_w2;
	wire_w_lg_dataa_sign_dffe1_wo345w(0) <= NOT dataa_sign_dffe1_wo;
	wire_w_lg_datab_sign_dffe1_wo348w(0) <= NOT datab_sign_dffe1_wo;
	wire_w_lg_denormal_result_w572w(0) <= NOT denormal_result_w;
	wire_w_lg_exp_amb_mux_dffe15_wo316w(0) <= NOT exp_amb_mux_dffe15_wo;
	wire_w_lg_exp_amb_mux_w275w(0) <= NOT exp_amb_mux_w;
	wire_w_lg_force_infinity_w643w(0) <= NOT force_infinity_w;
	wire_w_lg_force_nan_w644w(0) <= NOT force_nan_w;
	wire_w_lg_force_zero_w642w(0) <= NOT force_zero_w;
	wire_w_lg_input_dataa_denormal_dffe11_wo233w(0) <= NOT input_dataa_denormal_dffe11_wo;
	wire_w_lg_input_dataa_infinite_dffe11_wo246w(0) <= NOT input_dataa_infinite_dffe11_wo;
	wire_w_lg_input_dataa_zero_dffe11_wo245w(0) <= NOT input_dataa_zero_dffe11_wo;
	wire_w_lg_input_datab_denormal_dffe11_wo252w(0) <= NOT input_datab_denormal_dffe11_wo;
	wire_w_lg_input_datab_infinite_dffe11_wo265w(0) <= NOT input_datab_infinite_dffe11_wo;
	wire_w_lg_input_datab_infinite_dffe15_wo339w(0) <= NOT input_datab_infinite_dffe15_wo;
	wire_w_lg_input_datab_zero_dffe11_wo264w(0) <= NOT input_datab_zero_dffe11_wo;
	wire_w_lg_man_res_is_not_zero_dffe4_wo641w(0) <= NOT man_res_is_not_zero_dffe4_wo;
	wire_w_lg_man_res_not_zero_dffe26_wo517w(0) <= NOT man_res_not_zero_dffe26_wo;
	wire_w_lg_need_complement_dffe22_wo387w(0) <= NOT need_complement_dffe22_wo;
	wire_w_lg_sticky_bit_dffe1_wo357w(0) <= NOT sticky_bit_dffe1_wo;
	wire_w_lg_w_exp_adjustment2_add_sub_w_range525w574w(0) <= NOT wire_w_exp_adjustment2_add_sub_w_range525w(0);
	wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w291w(0) <= NOT wire_w_exp_diff_abs_exceed_max_w_range289w(0);
	wire_w_lg_w_man_a_not_zero_w_range215w219w(0) <= NOT wire_w_man_a_not_zero_w_range215w(0);
	wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range401w404w(0) <= NOT wire_w_man_add_sub_res_mag_dffe27_wo_range401w(0);
	wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) <= NOT wire_w_man_add_sub_res_mag_dffe27_wo_range395w(0);
	wire_w_lg_w_man_add_sub_w_range386w389w(0) <= NOT wire_w_man_add_sub_w_range386w(0);
	wire_w_lg_w_man_b_not_zero_w_range218w225w(0) <= NOT wire_w_man_b_not_zero_w_range218w(0);
	wire_w_lg_w_man_res_rounding_add_sub_w_range599w600w(0) <= NOT wire_w_man_res_rounding_add_sub_w_range599w(0);
	loop117 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_force_zero_w648w651w652w(i) <= wire_w_lg_w_lg_force_zero_w648w651w(i) OR wire_w_lg_w_lg_w_lg_force_zero_w648w649w650w(i);
	END GENERATE loop117;
	loop118 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_force_zero_w648w660w661w(i) <= wire_w_lg_w_lg_force_zero_w648w660w(i) OR wire_w_lg_w_lg_w_lg_force_zero_w648w649w659w(i);
	END GENERATE loop118;
	loop119 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_force_infinity_w654w655w(i) <= wire_w_lg_force_infinity_w654w(i) OR wire_w_lg_w_lg_force_infinity_w643w653w(i);
	END GENERATE loop119;
	loop120 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_force_infinity_w663w664w(i) <= wire_w_lg_force_infinity_w663w(i) OR wire_w_lg_w_lg_force_infinity_w643w662w(i);
	END GENERATE loop120;
	wire_w_lg_force_zero_w648w(0) <= force_zero_w OR denormal_flag_w;
	wire_w_lg_sticky_bit_dffe27_wo416w(0) <= sticky_bit_dffe27_wo OR wire_w_man_add_sub_res_mag_dffe27_wo_range410w(0);
	wire_w_lg_w_dataa_range141w142w(0) <= wire_w_dataa_range141w(0) OR wire_w_man_a_not_zero_w_range137w(0);
	wire_w_lg_w_dataa_range147w148w(0) <= wire_w_dataa_range147w(0) OR wire_w_man_a_not_zero_w_range143w(0);
	wire_w_lg_w_dataa_range153w154w(0) <= wire_w_dataa_range153w(0) OR wire_w_man_a_not_zero_w_range149w(0);
	wire_w_lg_w_dataa_range159w160w(0) <= wire_w_dataa_range159w(0) OR wire_w_man_a_not_zero_w_range155w(0);
	wire_w_lg_w_dataa_range165w166w(0) <= wire_w_dataa_range165w(0) OR wire_w_man_a_not_zero_w_range161w(0);
	wire_w_lg_w_dataa_range171w172w(0) <= wire_w_dataa_range171w(0) OR wire_w_man_a_not_zero_w_range167w(0);
	wire_w_lg_w_dataa_range177w178w(0) <= wire_w_dataa_range177w(0) OR wire_w_man_a_not_zero_w_range173w(0);
	wire_w_lg_w_dataa_range183w184w(0) <= wire_w_dataa_range183w(0) OR wire_w_man_a_not_zero_w_range179w(0);
	wire_w_lg_w_dataa_range189w190w(0) <= wire_w_dataa_range189w(0) OR wire_w_man_a_not_zero_w_range185w(0);
	wire_w_lg_w_dataa_range195w196w(0) <= wire_w_dataa_range195w(0) OR wire_w_man_a_not_zero_w_range191w(0);
	wire_w_lg_w_dataa_range87w88w(0) <= wire_w_dataa_range87w(0) OR wire_w_man_a_not_zero_w_range12w(0);
	wire_w_lg_w_dataa_range201w202w(0) <= wire_w_dataa_range201w(0) OR wire_w_man_a_not_zero_w_range197w(0);
	wire_w_lg_w_dataa_range207w208w(0) <= wire_w_dataa_range207w(0) OR wire_w_man_a_not_zero_w_range203w(0);
	wire_w_lg_w_dataa_range213w214w(0) <= wire_w_dataa_range213w(0) OR wire_w_man_a_not_zero_w_range209w(0);
	wire_w_lg_w_dataa_range17w18w(0) <= wire_w_dataa_range17w(0) OR wire_w_exp_a_not_zero_w_range2w(0);
	wire_w_lg_w_dataa_range27w28w(0) <= wire_w_dataa_range27w(0) OR wire_w_exp_a_not_zero_w_range19w(0);
	wire_w_lg_w_dataa_range37w38w(0) <= wire_w_dataa_range37w(0) OR wire_w_exp_a_not_zero_w_range29w(0);
	wire_w_lg_w_dataa_range47w48w(0) <= wire_w_dataa_range47w(0) OR wire_w_exp_a_not_zero_w_range39w(0);
	wire_w_lg_w_dataa_range57w58w(0) <= wire_w_dataa_range57w(0) OR wire_w_exp_a_not_zero_w_range49w(0);
	wire_w_lg_w_dataa_range67w68w(0) <= wire_w_dataa_range67w(0) OR wire_w_exp_a_not_zero_w_range59w(0);
	wire_w_lg_w_dataa_range93w94w(0) <= wire_w_dataa_range93w(0) OR wire_w_man_a_not_zero_w_range89w(0);
	wire_w_lg_w_dataa_range77w78w(0) <= wire_w_dataa_range77w(0) OR wire_w_exp_a_not_zero_w_range69w(0);
	wire_w_lg_w_dataa_range99w100w(0) <= wire_w_dataa_range99w(0) OR wire_w_man_a_not_zero_w_range95w(0);
	wire_w_lg_w_dataa_range105w106w(0) <= wire_w_dataa_range105w(0) OR wire_w_man_a_not_zero_w_range101w(0);
	wire_w_lg_w_dataa_range111w112w(0) <= wire_w_dataa_range111w(0) OR wire_w_man_a_not_zero_w_range107w(0);
	wire_w_lg_w_dataa_range117w118w(0) <= wire_w_dataa_range117w(0) OR wire_w_man_a_not_zero_w_range113w(0);
	wire_w_lg_w_dataa_range123w124w(0) <= wire_w_dataa_range123w(0) OR wire_w_man_a_not_zero_w_range119w(0);
	wire_w_lg_w_dataa_range129w130w(0) <= wire_w_dataa_range129w(0) OR wire_w_man_a_not_zero_w_range125w(0);
	wire_w_lg_w_dataa_range135w136w(0) <= wire_w_dataa_range135w(0) OR wire_w_man_a_not_zero_w_range131w(0);
	wire_w_lg_w_datab_range144w145w(0) <= wire_w_datab_range144w(0) OR wire_w_man_b_not_zero_w_range140w(0);
	wire_w_lg_w_datab_range150w151w(0) <= wire_w_datab_range150w(0) OR wire_w_man_b_not_zero_w_range146w(0);
	wire_w_lg_w_datab_range156w157w(0) <= wire_w_datab_range156w(0) OR wire_w_man_b_not_zero_w_range152w(0);
	wire_w_lg_w_datab_range162w163w(0) <= wire_w_datab_range162w(0) OR wire_w_man_b_not_zero_w_range158w(0);
	wire_w_lg_w_datab_range168w169w(0) <= wire_w_datab_range168w(0) OR wire_w_man_b_not_zero_w_range164w(0);
	wire_w_lg_w_datab_range174w175w(0) <= wire_w_datab_range174w(0) OR wire_w_man_b_not_zero_w_range170w(0);
	wire_w_lg_w_datab_range180w181w(0) <= wire_w_datab_range180w(0) OR wire_w_man_b_not_zero_w_range176w(0);
	wire_w_lg_w_datab_range186w187w(0) <= wire_w_datab_range186w(0) OR wire_w_man_b_not_zero_w_range182w(0);
	wire_w_lg_w_datab_range192w193w(0) <= wire_w_datab_range192w(0) OR wire_w_man_b_not_zero_w_range188w(0);
	wire_w_lg_w_datab_range198w199w(0) <= wire_w_datab_range198w(0) OR wire_w_man_b_not_zero_w_range194w(0);
	wire_w_lg_w_datab_range90w91w(0) <= wire_w_datab_range90w(0) OR wire_w_man_b_not_zero_w_range15w(0);
	wire_w_lg_w_datab_range204w205w(0) <= wire_w_datab_range204w(0) OR wire_w_man_b_not_zero_w_range200w(0);
	wire_w_lg_w_datab_range210w211w(0) <= wire_w_datab_range210w(0) OR wire_w_man_b_not_zero_w_range206w(0);
	wire_w_lg_w_datab_range216w217w(0) <= wire_w_datab_range216w(0) OR wire_w_man_b_not_zero_w_range212w(0);
	wire_w_lg_w_datab_range20w21w(0) <= wire_w_datab_range20w(0) OR wire_w_exp_b_not_zero_w_range5w(0);
	wire_w_lg_w_datab_range30w31w(0) <= wire_w_datab_range30w(0) OR wire_w_exp_b_not_zero_w_range22w(0);
	wire_w_lg_w_datab_range40w41w(0) <= wire_w_datab_range40w(0) OR wire_w_exp_b_not_zero_w_range32w(0);
	wire_w_lg_w_datab_range50w51w(0) <= wire_w_datab_range50w(0) OR wire_w_exp_b_not_zero_w_range42w(0);
	wire_w_lg_w_datab_range60w61w(0) <= wire_w_datab_range60w(0) OR wire_w_exp_b_not_zero_w_range52w(0);
	wire_w_lg_w_datab_range70w71w(0) <= wire_w_datab_range70w(0) OR wire_w_exp_b_not_zero_w_range62w(0);
	wire_w_lg_w_datab_range96w97w(0) <= wire_w_datab_range96w(0) OR wire_w_man_b_not_zero_w_range92w(0);
	wire_w_lg_w_datab_range80w81w(0) <= wire_w_datab_range80w(0) OR wire_w_exp_b_not_zero_w_range72w(0);
	wire_w_lg_w_datab_range102w103w(0) <= wire_w_datab_range102w(0) OR wire_w_man_b_not_zero_w_range98w(0);
	wire_w_lg_w_datab_range108w109w(0) <= wire_w_datab_range108w(0) OR wire_w_man_b_not_zero_w_range104w(0);
	wire_w_lg_w_datab_range114w115w(0) <= wire_w_datab_range114w(0) OR wire_w_man_b_not_zero_w_range110w(0);
	wire_w_lg_w_datab_range120w121w(0) <= wire_w_datab_range120w(0) OR wire_w_man_b_not_zero_w_range116w(0);
	wire_w_lg_w_datab_range126w127w(0) <= wire_w_datab_range126w(0) OR wire_w_man_b_not_zero_w_range122w(0);
	wire_w_lg_w_datab_range132w133w(0) <= wire_w_datab_range132w(0) OR wire_w_man_b_not_zero_w_range128w(0);
	wire_w_lg_w_datab_range138w139w(0) <= wire_w_datab_range138w(0) OR wire_w_man_b_not_zero_w_range134w(0);
	wire_w_lg_w_exp_diff_abs_exceed_max_w_range282w285w(0) <= wire_w_exp_diff_abs_exceed_max_w_range282w(0) OR wire_w_exp_diff_abs_w_range284w(0);
	wire_w_lg_w_exp_diff_abs_exceed_max_w_range286w288w(0) <= wire_w_exp_diff_abs_exceed_max_w_range286w(0) OR wire_w_exp_diff_abs_w_range287w(0);
	wire_w_lg_w_exp_res_not_zero_w_range530w533w(0) <= wire_w_exp_res_not_zero_w_range530w(0) OR wire_w_exp_adjustment2_add_sub_w_range532w(0);
	wire_w_lg_w_exp_res_not_zero_w_range534w536w(0) <= wire_w_exp_res_not_zero_w_range534w(0) OR wire_w_exp_adjustment2_add_sub_w_range535w(0);
	wire_w_lg_w_exp_res_not_zero_w_range537w539w(0) <= wire_w_exp_res_not_zero_w_range537w(0) OR wire_w_exp_adjustment2_add_sub_w_range538w(0);
	wire_w_lg_w_exp_res_not_zero_w_range540w542w(0) <= wire_w_exp_res_not_zero_w_range540w(0) OR wire_w_exp_adjustment2_add_sub_w_range541w(0);
	wire_w_lg_w_exp_res_not_zero_w_range543w545w(0) <= wire_w_exp_res_not_zero_w_range543w(0) OR wire_w_exp_adjustment2_add_sub_w_range544w(0);
	wire_w_lg_w_exp_res_not_zero_w_range546w548w(0) <= wire_w_exp_res_not_zero_w_range546w(0) OR wire_w_exp_adjustment2_add_sub_w_range547w(0);
	wire_w_lg_w_exp_res_not_zero_w_range549w551w(0) <= wire_w_exp_res_not_zero_w_range549w(0) OR wire_w_exp_adjustment2_add_sub_w_range550w(0);
	wire_w_lg_w_exp_res_not_zero_w_range552w553w(0) <= wire_w_exp_res_not_zero_w_range552w(0) OR wire_w_exp_adjustment2_add_sub_w_range525w(0);
	wire_w_lg_w_man_res_not_zero_w2_range431w434w(0) <= wire_w_man_res_not_zero_w2_range431w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range433w(0);
	wire_w_lg_w_man_res_not_zero_w2_range462w464w(0) <= wire_w_man_res_not_zero_w2_range462w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range463w(0);
	wire_w_lg_w_man_res_not_zero_w2_range465w467w(0) <= wire_w_man_res_not_zero_w2_range465w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range466w(0);
	wire_w_lg_w_man_res_not_zero_w2_range468w470w(0) <= wire_w_man_res_not_zero_w2_range468w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range469w(0);
	wire_w_lg_w_man_res_not_zero_w2_range471w473w(0) <= wire_w_man_res_not_zero_w2_range471w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range472w(0);
	wire_w_lg_w_man_res_not_zero_w2_range474w476w(0) <= wire_w_man_res_not_zero_w2_range474w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range475w(0);
	wire_w_lg_w_man_res_not_zero_w2_range477w479w(0) <= wire_w_man_res_not_zero_w2_range477w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range478w(0);
	wire_w_lg_w_man_res_not_zero_w2_range480w482w(0) <= wire_w_man_res_not_zero_w2_range480w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range481w(0);
	wire_w_lg_w_man_res_not_zero_w2_range483w485w(0) <= wire_w_man_res_not_zero_w2_range483w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range484w(0);
	wire_w_lg_w_man_res_not_zero_w2_range486w488w(0) <= wire_w_man_res_not_zero_w2_range486w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range487w(0);
	wire_w_lg_w_man_res_not_zero_w2_range489w491w(0) <= wire_w_man_res_not_zero_w2_range489w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range490w(0);
	wire_w_lg_w_man_res_not_zero_w2_range435w437w(0) <= wire_w_man_res_not_zero_w2_range435w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range436w(0);
	wire_w_lg_w_man_res_not_zero_w2_range492w494w(0) <= wire_w_man_res_not_zero_w2_range492w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range493w(0);
	wire_w_lg_w_man_res_not_zero_w2_range495w497w(0) <= wire_w_man_res_not_zero_w2_range495w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range496w(0);
	wire_w_lg_w_man_res_not_zero_w2_range498w500w(0) <= wire_w_man_res_not_zero_w2_range498w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range499w(0);
	wire_w_lg_w_man_res_not_zero_w2_range501w503w(0) <= wire_w_man_res_not_zero_w2_range501w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range502w(0);
	wire_w_lg_w_man_res_not_zero_w2_range438w440w(0) <= wire_w_man_res_not_zero_w2_range438w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range439w(0);
	wire_w_lg_w_man_res_not_zero_w2_range441w443w(0) <= wire_w_man_res_not_zero_w2_range441w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range442w(0);
	wire_w_lg_w_man_res_not_zero_w2_range444w446w(0) <= wire_w_man_res_not_zero_w2_range444w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range445w(0);
	wire_w_lg_w_man_res_not_zero_w2_range447w449w(0) <= wire_w_man_res_not_zero_w2_range447w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range448w(0);
	wire_w_lg_w_man_res_not_zero_w2_range450w452w(0) <= wire_w_man_res_not_zero_w2_range450w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range451w(0);
	wire_w_lg_w_man_res_not_zero_w2_range453w455w(0) <= wire_w_man_res_not_zero_w2_range453w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range454w(0);
	wire_w_lg_w_man_res_not_zero_w2_range456w458w(0) <= wire_w_man_res_not_zero_w2_range456w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range457w(0);
	wire_w_lg_w_man_res_not_zero_w2_range459w461w(0) <= wire_w_man_res_not_zero_w2_range459w(0) OR wire_w_man_add_sub_res_mag_dffe21_wo_range460w(0);
	wire_w_lg_aligned_datab_sign_dffe15_wo336w(0) <= aligned_datab_sign_dffe15_wo XOR add_sub_dffe15_wo;
	aclr <= '0';
	add_sub_dffe11_wi <= add_sub;
	add_sub_dffe11_wo <= add_sub_dffe11_wi;
	add_sub_dffe12_wi <= add_sub_dffe11_wo;
	add_sub_dffe12_wo <= add_sub_dffe12_wi;
	add_sub_dffe13_wi <= add_sub_dffe12_wo;
	add_sub_dffe13_wo <= add_sub_dffe13_wi;
	add_sub_dffe14_wi <= add_sub_dffe13_wo;
	add_sub_dffe14_wo <= add_sub_dffe14_wi;
	add_sub_dffe15_wi <= add_sub_dffe14_wo;
	add_sub_dffe15_wo <= add_sub_dffe15_wi;
	add_sub_dffe1_wi <= add_sub_dffe15_wo;
	add_sub_dffe1_wo <= add_sub_dffe1;
	add_sub_dffe25_wi <= add_sub_w2;
	add_sub_dffe25_wo <= add_sub_dffe25_wi;
	add_sub_w2 <= ((((wire_w_lg_dataa_sign_dffe1_wo351w(0) AND wire_w_lg_add_sub_dffe1_wo344w(0)) OR wire_w_lg_w_lg_w_lg_dataa_sign_dffe1_wo345w349w350w(0)) OR (wire_w_lg_w_lg_dataa_sign_dffe1_wo345w346w(0) AND wire_w_lg_add_sub_dffe1_wo344w(0))) OR wire_w_lg_w_lg_dataa_sign_dffe1_wo342w343w(0));
	adder_upper_w <= man_intermediate_res_w(25 DOWNTO 13);
	aligned_dataa_exp_dffe12_wi <= aligned_dataa_exp_w;
	aligned_dataa_exp_dffe12_wo <= aligned_dataa_exp_dffe12_wi;
	aligned_dataa_exp_dffe13_wi <= aligned_dataa_exp_dffe12_wo;
	aligned_dataa_exp_dffe13_wo <= aligned_dataa_exp_dffe13_wi;
	aligned_dataa_exp_dffe14_wi <= aligned_dataa_exp_dffe13_wo;
	aligned_dataa_exp_dffe14_wo <= aligned_dataa_exp_dffe14_wi;
	aligned_dataa_exp_dffe15_wi <= aligned_dataa_exp_dffe14_wo;
	aligned_dataa_exp_dffe15_wo <= aligned_dataa_exp_dffe15_wi;
	aligned_dataa_exp_w <= ( "0" & wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w234w);
	aligned_dataa_man_dffe12_wi <= aligned_dataa_man_w(25 DOWNTO 2);
	aligned_dataa_man_dffe12_wo <= aligned_dataa_man_dffe12_wi;
	aligned_dataa_man_dffe13_wi <= aligned_dataa_man_dffe12_wo;
	aligned_dataa_man_dffe13_wo <= aligned_dataa_man_dffe13_wi;
	aligned_dataa_man_dffe14_wi <= aligned_dataa_man_dffe13_wo;
	aligned_dataa_man_dffe14_wo <= aligned_dataa_man_dffe14_wi;
	aligned_dataa_man_dffe15_w <= ( aligned_dataa_man_dffe15_wo & "00");
	aligned_dataa_man_dffe15_wi <= aligned_dataa_man_dffe14_wo;
	aligned_dataa_man_dffe15_wo <= aligned_dataa_man_dffe15_wi;
	aligned_dataa_man_w <= ( wire_w248w & wire_w_lg_w_lg_input_dataa_denormal_dffe11_wo233w243w & "00");
	aligned_dataa_sign_dffe12_wi <= aligned_dataa_sign_w;
	aligned_dataa_sign_dffe12_wo <= aligned_dataa_sign_dffe12_wi;
	aligned_dataa_sign_dffe13_wi <= aligned_dataa_sign_dffe12_wo;
	aligned_dataa_sign_dffe13_wo <= aligned_dataa_sign_dffe13_wi;
	aligned_dataa_sign_dffe14_wi <= aligned_dataa_sign_dffe13_wo;
	aligned_dataa_sign_dffe14_wo <= aligned_dataa_sign_dffe14_wi;
	aligned_dataa_sign_dffe15_wi <= aligned_dataa_sign_dffe14_wo;
	aligned_dataa_sign_dffe15_wo <= aligned_dataa_sign_dffe15_wi;
	aligned_dataa_sign_w <= dataa_dffe11_wo(31);
	aligned_datab_exp_dffe12_wi <= aligned_datab_exp_w;
	aligned_datab_exp_dffe12_wo <= aligned_datab_exp_dffe12_wi;
	aligned_datab_exp_dffe13_wi <= aligned_datab_exp_dffe12_wo;
	aligned_datab_exp_dffe13_wo <= aligned_datab_exp_dffe13_wi;
	aligned_datab_exp_dffe14_wi <= aligned_datab_exp_dffe13_wo;
	aligned_datab_exp_dffe14_wo <= aligned_datab_exp_dffe14_wi;
	aligned_datab_exp_dffe15_wi <= aligned_datab_exp_dffe14_wo;
	aligned_datab_exp_dffe15_wo <= aligned_datab_exp_dffe15_wi;
	aligned_datab_exp_w <= ( "0" & wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w253w);
	aligned_datab_man_dffe12_wi <= aligned_datab_man_w(25 DOWNTO 2);
	aligned_datab_man_dffe12_wo <= aligned_datab_man_dffe12_wi;
	aligned_datab_man_dffe13_wi <= aligned_datab_man_dffe12_wo;
	aligned_datab_man_dffe13_wo <= aligned_datab_man_dffe13_wi;
	aligned_datab_man_dffe14_wi <= aligned_datab_man_dffe13_wo;
	aligned_datab_man_dffe14_wo <= aligned_datab_man_dffe14_wi;
	aligned_datab_man_dffe15_w <= ( aligned_datab_man_dffe15_wo & "00");
	aligned_datab_man_dffe15_wi <= aligned_datab_man_dffe14_wo;
	aligned_datab_man_dffe15_wo <= aligned_datab_man_dffe15_wi;
	aligned_datab_man_w <= ( wire_w267w & wire_w_lg_w_lg_input_datab_denormal_dffe11_wo252w262w & "00");
	aligned_datab_sign_dffe12_wi <= aligned_datab_sign_w;
	aligned_datab_sign_dffe12_wo <= aligned_datab_sign_dffe12_wi;
	aligned_datab_sign_dffe13_wi <= aligned_datab_sign_dffe12_wo;
	aligned_datab_sign_dffe13_wo <= aligned_datab_sign_dffe13_wi;
	aligned_datab_sign_dffe14_wi <= aligned_datab_sign_dffe13_wo;
	aligned_datab_sign_dffe14_wo <= aligned_datab_sign_dffe14_wi;
	aligned_datab_sign_dffe15_wi <= aligned_datab_sign_dffe14_wo;
	aligned_datab_sign_dffe15_wo <= aligned_datab_sign_dffe15_wi;
	aligned_datab_sign_w <= datab_dffe11_wo(31);
	borrow_w <= (wire_w_lg_sticky_bit_dffe1_wo357w(0) AND wire_w_lg_add_sub_w2356w(0));
	both_inputs_are_infinite_dffe1_wi <= (input_dataa_infinite_dffe15_wo AND input_datab_infinite_dffe15_wo);
	both_inputs_are_infinite_dffe1_wo <= both_inputs_are_infinite_dffe1;
	both_inputs_are_infinite_dffe25_wi <= both_inputs_are_infinite_dffe1_wo;
	both_inputs_are_infinite_dffe25_wo <= both_inputs_are_infinite_dffe25_wi;
	clk_en <= '1';
	data_exp_dffe1_wi <= (wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w317w OR wire_w_lg_exp_amb_mux_dffe15_wo314w);
	data_exp_dffe1_wo <= data_exp_dffe1;
	dataa_dffe11_wi <= dataa;
	dataa_dffe11_wo <= dataa_dffe11_wi;
	dataa_man_dffe1_wi <= (wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w324w OR wire_w_lg_exp_amb_mux_dffe15_wo323w);
	dataa_man_dffe1_wo <= dataa_man_dffe1;
	dataa_sign_dffe1_wi <= aligned_dataa_sign_dffe15_wo;
	dataa_sign_dffe1_wo <= dataa_sign_dffe1;
	dataa_sign_dffe25_wi <= dataa_sign_dffe1_wo;
	dataa_sign_dffe25_wo <= dataa_sign_dffe25_wi;
	datab_dffe11_wi <= datab;
	datab_dffe11_wo <= datab_dffe11_wi;
	datab_man_dffe1_wi <= (wire_w_lg_w_lg_exp_amb_mux_dffe15_wo316w331w OR wire_w_lg_exp_amb_mux_dffe15_wo330w);
	datab_man_dffe1_wo <= datab_man_dffe1;
	datab_sign_dffe1_wi <= aligned_datab_sign_dffe15_wo;
	datab_sign_dffe1_wo <= datab_sign_dffe1;
	denormal_flag_w <= (((wire_w_lg_force_nan_w644w(0) AND wire_w_lg_force_infinity_w643w(0)) AND wire_w_lg_force_zero_w642w(0)) AND denormal_res_dffe4_wo);
	denormal_res_dffe32_wi <= denormal_result_w;
	denormal_res_dffe32_wo <= denormal_res_dffe32_wi;
	denormal_res_dffe33_wi <= denormal_res_dffe32_wo;
	denormal_res_dffe33_wo <= denormal_res_dffe33_wi;
	denormal_res_dffe3_wi <= denormal_res_dffe33_wo;
	denormal_res_dffe3_wo <= denormal_res_dffe3;
	denormal_res_dffe41_wi <= denormal_res_dffe42_wo;
	denormal_res_dffe41_wo <= denormal_res_dffe41_wi;
	denormal_res_dffe42_wi <= denormal_res_dffe3_wo;
	denormal_res_dffe42_wo <= denormal_res_dffe42_wi;
	denormal_res_dffe4_wi <= denormal_res_dffe41_wo;
	denormal_res_dffe4_wo <= denormal_res_dffe4;
	denormal_result_w <= ((NOT exp_res_not_zero_w(8)) OR exp_adjustment2_add_sub_w(8));
	exp_a_all_one_w <= ( wire_w_lg_w_dataa_range77w83w & wire_w_lg_w_dataa_range67w73w & wire_w_lg_w_dataa_range57w63w & wire_w_lg_w_dataa_range47w53w & wire_w_lg_w_dataa_range37w43w & wire_w_lg_w_dataa_range27w33w & wire_w_lg_w_dataa_range17w23w & dataa(23));
	exp_a_not_zero_w <= ( wire_w_lg_w_dataa_range77w78w & wire_w_lg_w_dataa_range67w68w & wire_w_lg_w_dataa_range57w58w & wire_w_lg_w_dataa_range47w48w & wire_w_lg_w_dataa_range37w38w & wire_w_lg_w_dataa_range27w28w & wire_w_lg_w_dataa_range17w18w & dataa(23));
	exp_adj_0pads <= (OTHERS => '0');
	exp_adj_dffe21_wi <= (wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w398w OR wire_w397w);
	exp_adj_dffe21_wo <= exp_adj_dffe21;
	exp_adj_dffe23_wi <= exp_adj_dffe21_wo;
	exp_adj_dffe23_wo <= exp_adj_dffe23_wi;
	exp_adj_dffe26_wi <= exp_adj_dffe23_wo;
	exp_adj_dffe26_wo <= exp_adj_dffe26_wi;
	exp_adjust_by_add1 <= "01";
	exp_adjust_by_add2 <= "10";
	exp_adjustment2_add_sub_dataa_w <= exp_value;
	exp_adjustment2_add_sub_datab_w <= exp_adjustment_add_sub_w;
	exp_adjustment2_add_sub_w <= wire_add_sub5_result;
	exp_adjustment_add_sub_dataa_w <= ( priority_encoder_1pads_w & wire_leading_zeroes_cnt_q);
	exp_adjustment_add_sub_datab_w <= ( exp_adj_0pads & exp_adj_dffe26_wo);
	exp_adjustment_add_sub_w <= wire_add_sub4_result;
	exp_all_ones_w <= (OTHERS => '1');
	exp_all_zeros_w <= (OTHERS => '0');
	exp_amb_mux_dffe13_wi <= exp_amb_mux_w;
	exp_amb_mux_dffe13_wo <= exp_amb_mux_dffe13_wi;
	exp_amb_mux_dffe14_wi <= exp_amb_mux_dffe13_wo;
	exp_amb_mux_dffe14_wo <= exp_amb_mux_dffe14_wi;
	exp_amb_mux_dffe15_wi <= exp_amb_mux_dffe14_wo;
	exp_amb_mux_dffe15_wo <= exp_amb_mux_dffe15_wi;
	exp_amb_mux_w <= exp_amb_w(8);
	exp_amb_w <= wire_add_sub1_result;
	exp_b_all_one_w <= ( wire_w_lg_w_datab_range80w85w & wire_w_lg_w_datab_range70w75w & wire_w_lg_w_datab_range60w65w & wire_w_lg_w_datab_range50w55w & wire_w_lg_w_datab_range40w45w & wire_w_lg_w_datab_range30w35w & wire_w_lg_w_datab_range20w25w & datab(23));
	exp_b_not_zero_w <= ( wire_w_lg_w_datab_range80w81w & wire_w_lg_w_datab_range70w71w & wire_w_lg_w_datab_range60w61w & wire_w_lg_w_datab_range50w51w & wire_w_lg_w_datab_range40w41w & wire_w_lg_w_datab_range30w31w & wire_w_lg_w_datab_range20w21w & datab(23));
	exp_bma_w <= wire_add_sub2_result;
	exp_diff_abs_exceed_max_w <= ( wire_w_lg_w_exp_diff_abs_exceed_max_w_range286w288w & wire_w_lg_w_exp_diff_abs_exceed_max_w_range282w285w & exp_diff_abs_w(5));
	exp_diff_abs_max_w <= (OTHERS => '1');
	exp_diff_abs_w <= (wire_w_lg_w_lg_exp_amb_mux_w275w276w OR wire_w_lg_exp_amb_mux_w273w);
	exp_intermediate_res_dffe41_wi <= exp_intermediate_res_dffe42_wo;
	exp_intermediate_res_dffe41_wo <= exp_intermediate_res_dffe41_wi;
	exp_intermediate_res_dffe42_wi <= exp_intermediate_res_w;
	exp_intermediate_res_dffe42_wo <= exp_intermediate_res_dffe42_wi;
	exp_intermediate_res_w <= exp_res_dffe3_wo;
	exp_out_dffe5_wi <= (wire_w_lg_force_nan_w657w OR wire_w_lg_w_lg_force_nan_w644w656w);
	exp_out_dffe5_wo <= exp_out_dffe5;
	exp_res_dffe21_wi <= exp_res_dffe27_wo;
	exp_res_dffe21_wo <= exp_res_dffe21;
	exp_res_dffe22_wi <= exp_res_dffe2_wo;
	exp_res_dffe22_wo <= exp_res_dffe22_wi;
	exp_res_dffe23_wi <= exp_res_dffe21_wo;
	exp_res_dffe23_wo <= exp_res_dffe23_wi;
	exp_res_dffe25_wi <= data_exp_dffe1_wo;
	exp_res_dffe25_wo <= exp_res_dffe25_wi;
	exp_res_dffe26_wi <= exp_res_dffe23_wo;
	exp_res_dffe26_wo <= exp_res_dffe26_wi;
	exp_res_dffe27_wi <= exp_res_dffe22_wo;
	exp_res_dffe27_wo <= exp_res_dffe27_wi;
	exp_res_dffe2_wi <= exp_res_dffe25_wo;
	exp_res_dffe2_wo <= exp_res_dffe2;
	exp_res_dffe32_wi <= wire_w_lg_w_lg_denormal_result_w572w573w;
	exp_res_dffe32_wo <= exp_res_dffe32_wi;
	exp_res_dffe33_wi <= exp_res_dffe32_wo;
	exp_res_dffe33_wo <= exp_res_dffe33_wi;
	exp_res_dffe3_wi <= exp_res_dffe33_wo;
	exp_res_dffe3_wo <= exp_res_dffe3;
	exp_res_dffe4_wi <= exp_rounded_res_w;
	exp_res_dffe4_wo <= exp_res_dffe4;
	exp_res_max_w <= ( wire_w_lg_w_exp_res_max_w_range567w568w & wire_w_lg_w_exp_res_max_w_range565w566w & wire_w_lg_w_exp_res_max_w_range563w564w & wire_w_lg_w_exp_res_max_w_range561w562w & wire_w_lg_w_exp_res_max_w_range559w560w & wire_w_lg_w_exp_res_max_w_range557w558w & wire_w_lg_w_exp_res_max_w_range554w556w & exp_adjustment2_add_sub_w(0));
	exp_res_not_zero_w <= ( wire_w_lg_w_exp_res_not_zero_w_range552w553w & wire_w_lg_w_exp_res_not_zero_w_range549w551w & wire_w_lg_w_exp_res_not_zero_w_range546w548w & wire_w_lg_w_exp_res_not_zero_w_range543w545w & wire_w_lg_w_exp_res_not_zero_w_range540w542w & wire_w_lg_w_exp_res_not_zero_w_range537w539w & wire_w_lg_w_exp_res_not_zero_w_range534w536w & wire_w_lg_w_exp_res_not_zero_w_range530w533w & exp_adjustment2_add_sub_w(0));
	exp_res_rounding_adder_dataa_w <= ( "0" & exp_intermediate_res_dffe41_wo);
	exp_res_rounding_adder_w <= wire_add_sub6_result;
	exp_rounded_res_infinity_w <= exp_rounded_res_max_w(7);
	exp_rounded_res_max_w <= ( wire_w_lg_w_exp_rounded_res_max_w_range634w636w & wire_w_lg_w_exp_rounded_res_max_w_range631w633w & wire_w_lg_w_exp_rounded_res_max_w_range628w630w & wire_w_lg_w_exp_rounded_res_max_w_range625w627w & wire_w_lg_w_exp_rounded_res_max_w_range622w624w & wire_w_lg_w_exp_rounded_res_max_w_range619w621w & wire_w_lg_w_exp_rounded_res_max_w_range615w618w & exp_rounded_res_w(0));
	exp_rounded_res_w <= exp_res_rounding_adder_w(7 DOWNTO 0);
	exp_rounding_adjustment_w <= ( "00000000" & man_res_rounding_add_sub_w(24));
	exp_value <= ( "0" & exp_res_dffe26_wo);
	force_infinity_w <= ((input_is_infinite_dffe4_wo OR rounded_res_infinity_dffe4_wo) OR infinite_res_dffe4_wo);
	force_nan_w <= (infinity_magnitude_sub_dffe4_wo OR input_is_nan_dffe4_wo);
	force_zero_w <= wire_w_lg_man_res_is_not_zero_dffe4_wo641w(0);
	guard_bit_dffe3_wo <= man_res_w3(0);
	infinite_output_sign_dffe1_wi <= (wire_w_lg_w_lg_input_datab_infinite_dffe15_wo339w340w(0) OR wire_w_lg_input_datab_infinite_dffe15_wo338w(0));
	infinite_output_sign_dffe1_wo <= infinite_output_sign_dffe1;
	infinite_output_sign_dffe21_wi <= infinite_output_sign_dffe27_wo;
	infinite_output_sign_dffe21_wo <= infinite_output_sign_dffe21;
	infinite_output_sign_dffe22_wi <= infinite_output_sign_dffe2_wo;
	infinite_output_sign_dffe22_wo <= infinite_output_sign_dffe22_wi;
	infinite_output_sign_dffe23_wi <= infinite_output_sign_dffe21_wo;
	infinite_output_sign_dffe23_wo <= infinite_output_sign_dffe23_wi;
	infinite_output_sign_dffe25_wi <= infinite_output_sign_dffe1_wo;
	infinite_output_sign_dffe25_wo <= infinite_output_sign_dffe25_wi;
	infinite_output_sign_dffe26_wi <= infinite_output_sign_dffe23_wo;
	infinite_output_sign_dffe26_wo <= infinite_output_sign_dffe26_wi;
	infinite_output_sign_dffe27_wi <= infinite_output_sign_dffe22_wo;
	infinite_output_sign_dffe27_wo <= infinite_output_sign_dffe27_wi;
	infinite_output_sign_dffe2_wi <= infinite_output_sign_dffe25_wo;
	infinite_output_sign_dffe2_wo <= infinite_output_sign_dffe2;
	infinite_output_sign_dffe31_wi <= infinite_output_sign_dffe26_wo;
	infinite_output_sign_dffe31_wo <= infinite_output_sign_dffe31;
	infinite_output_sign_dffe32_wi <= infinite_output_sign_dffe31_wo;
	infinite_output_sign_dffe32_wo <= infinite_output_sign_dffe32_wi;
	infinite_output_sign_dffe33_wi <= infinite_output_sign_dffe32_wo;
	infinite_output_sign_dffe33_wo <= infinite_output_sign_dffe33_wi;
	infinite_output_sign_dffe3_wi <= infinite_output_sign_dffe33_wo;
	infinite_output_sign_dffe3_wo <= infinite_output_sign_dffe3;
	infinite_output_sign_dffe41_wi <= infinite_output_sign_dffe42_wo;
	infinite_output_sign_dffe41_wo <= infinite_output_sign_dffe41_wi;
	infinite_output_sign_dffe42_wi <= infinite_output_sign_dffe3_wo;
	infinite_output_sign_dffe42_wo <= infinite_output_sign_dffe42_wi;
	infinite_output_sign_dffe4_wi <= infinite_output_sign_dffe41_wo;
	infinite_output_sign_dffe4_wo <= infinite_output_sign_dffe4;
	infinite_res_dff32_wi <= wire_w_lg_w_exp_res_max_w_range569w575w(0);
	infinite_res_dff32_wo <= infinite_res_dff32_wi;
	infinite_res_dff33_wi <= infinite_res_dff32_wo;
	infinite_res_dff33_wo <= infinite_res_dff33_wi;
	infinite_res_dffe3_wi <= infinite_res_dff33_wo;
	infinite_res_dffe3_wo <= infinite_res_dffe3;
	infinite_res_dffe41_wi <= infinite_res_dffe42_wo;
	infinite_res_dffe41_wo <= infinite_res_dffe41_wi;
	infinite_res_dffe42_wi <= infinite_res_dffe3_wo;
	infinite_res_dffe42_wo <= infinite_res_dffe42_wi;
	infinite_res_dffe4_wi <= infinite_res_dffe41_wo;
	infinite_res_dffe4_wo <= infinite_res_dffe4;
	infinity_magnitude_sub_dffe21_wi <= infinity_magnitude_sub_dffe27_wo;
	infinity_magnitude_sub_dffe21_wo <= infinity_magnitude_sub_dffe21;
	infinity_magnitude_sub_dffe22_wi <= infinity_magnitude_sub_dffe2_wo;
	infinity_magnitude_sub_dffe22_wo <= infinity_magnitude_sub_dffe22_wi;
	infinity_magnitude_sub_dffe23_wi <= infinity_magnitude_sub_dffe21_wo;
	infinity_magnitude_sub_dffe23_wo <= infinity_magnitude_sub_dffe23_wi;
	infinity_magnitude_sub_dffe26_wi <= infinity_magnitude_sub_dffe23_wo;
	infinity_magnitude_sub_dffe26_wo <= infinity_magnitude_sub_dffe26_wi;
	infinity_magnitude_sub_dffe27_wi <= infinity_magnitude_sub_dffe22_wo;
	infinity_magnitude_sub_dffe27_wo <= infinity_magnitude_sub_dffe27_wi;
	infinity_magnitude_sub_dffe2_wi <= (wire_w_lg_add_sub_dffe25_wo505w(0) AND both_inputs_are_infinite_dffe25_wo);
	infinity_magnitude_sub_dffe2_wo <= infinity_magnitude_sub_dffe2;
	infinity_magnitude_sub_dffe31_wi <= infinity_magnitude_sub_dffe26_wo;
	infinity_magnitude_sub_dffe31_wo <= infinity_magnitude_sub_dffe31;
	infinity_magnitude_sub_dffe32_wi <= infinity_magnitude_sub_dffe31_wo;
	infinity_magnitude_sub_dffe32_wo <= infinity_magnitude_sub_dffe32_wi;
	infinity_magnitude_sub_dffe33_wi <= infinity_magnitude_sub_dffe32_wo;
	infinity_magnitude_sub_dffe33_wo <= infinity_magnitude_sub_dffe33_wi;
	infinity_magnitude_sub_dffe3_wi <= infinity_magnitude_sub_dffe33_wo;
	infinity_magnitude_sub_dffe3_wo <= infinity_magnitude_sub_dffe3;
	infinity_magnitude_sub_dffe41_wi <= infinity_magnitude_sub_dffe42_wo;
	infinity_magnitude_sub_dffe41_wo <= infinity_magnitude_sub_dffe41_wi;
	infinity_magnitude_sub_dffe42_wi <= infinity_magnitude_sub_dffe3_wo;
	infinity_magnitude_sub_dffe42_wo <= infinity_magnitude_sub_dffe42_wi;
	infinity_magnitude_sub_dffe4_wi <= infinity_magnitude_sub_dffe41_wo;
	infinity_magnitude_sub_dffe4_wo <= infinity_magnitude_sub_dffe4;
	input_dataa_denormal_dffe11_wi <= input_dataa_denormal_w;
	input_dataa_denormal_dffe11_wo <= input_dataa_denormal_dffe11_wi;
	input_dataa_denormal_w <= ((NOT exp_a_not_zero_w(7)) AND man_a_not_zero_w(22));
	input_dataa_infinite_dffe11_wi <= input_dataa_infinite_w;
	input_dataa_infinite_dffe11_wo <= input_dataa_infinite_dffe11_wi;
	input_dataa_infinite_dffe12_wi <= input_dataa_infinite_dffe11_wo;
	input_dataa_infinite_dffe12_wo <= input_dataa_infinite_dffe12_wi;
	input_dataa_infinite_dffe13_wi <= input_dataa_infinite_dffe12_wo;
	input_dataa_infinite_dffe13_wo <= input_dataa_infinite_dffe13_wi;
	input_dataa_infinite_dffe14_wi <= input_dataa_infinite_dffe13_wo;
	input_dataa_infinite_dffe14_wo <= input_dataa_infinite_dffe14_wi;
	input_dataa_infinite_dffe15_wi <= input_dataa_infinite_dffe14_wo;
	input_dataa_infinite_dffe15_wo <= input_dataa_infinite_dffe15_wi;
	input_dataa_infinite_w <= wire_w_lg_w_exp_a_all_one_w_range84w220w(0);
	input_dataa_nan_dffe11_wi <= input_dataa_nan_w;
	input_dataa_nan_dffe11_wo <= input_dataa_nan_dffe11_wi;
	input_dataa_nan_dffe12_wi <= input_dataa_nan_dffe11_wo;
	input_dataa_nan_dffe12_wo <= input_dataa_nan_dffe12_wi;
	input_dataa_nan_w <= (exp_a_all_one_w(7) AND man_a_not_zero_w(22));
	input_dataa_zero_dffe11_wi <= input_dataa_zero_w;
	input_dataa_zero_dffe11_wo <= input_dataa_zero_dffe11_wi;
	input_dataa_zero_w <= ((NOT exp_a_not_zero_w(7)) AND wire_w_lg_w_man_a_not_zero_w_range215w219w(0));
	input_datab_denormal_dffe11_wi <= input_datab_denormal_w;
	input_datab_denormal_dffe11_wo <= input_datab_denormal_dffe11_wi;
	input_datab_denormal_w <= ((NOT exp_b_not_zero_w(7)) AND man_b_not_zero_w(22));
	input_datab_infinite_dffe11_wi <= input_datab_infinite_w;
	input_datab_infinite_dffe11_wo <= input_datab_infinite_dffe11_wi;
	input_datab_infinite_dffe12_wi <= input_datab_infinite_dffe11_wo;
	input_datab_infinite_dffe12_wo <= input_datab_infinite_dffe12_wi;
	input_datab_infinite_dffe13_wi <= input_datab_infinite_dffe12_wo;
	input_datab_infinite_dffe13_wo <= input_datab_infinite_dffe13_wi;
	input_datab_infinite_dffe14_wi <= input_datab_infinite_dffe13_wo;
	input_datab_infinite_dffe14_wo <= input_datab_infinite_dffe14_wi;
	input_datab_infinite_dffe15_wi <= input_datab_infinite_dffe14_wo;
	input_datab_infinite_dffe15_wo <= input_datab_infinite_dffe15_wi;
	input_datab_infinite_w <= wire_w_lg_w_exp_b_all_one_w_range86w226w(0);
	input_datab_nan_dffe11_wi <= input_datab_nan_w;
	input_datab_nan_dffe11_wo <= input_datab_nan_dffe11_wi;
	input_datab_nan_dffe12_wi <= input_datab_nan_dffe11_wo;
	input_datab_nan_dffe12_wo <= input_datab_nan_dffe12_wi;
	input_datab_nan_w <= (exp_b_all_one_w(7) AND man_b_not_zero_w(22));
	input_datab_zero_dffe11_wi <= input_datab_zero_w;
	input_datab_zero_dffe11_wo <= input_datab_zero_dffe11_wi;
	input_datab_zero_w <= ((NOT exp_b_not_zero_w(7)) AND wire_w_lg_w_man_b_not_zero_w_range218w225w(0));
	input_is_infinite_dffe1_wi <= (input_dataa_infinite_dffe15_wo OR input_datab_infinite_dffe15_wo);
	input_is_infinite_dffe1_wo <= input_is_infinite_dffe1;
	input_is_infinite_dffe21_wi <= input_is_infinite_dffe27_wo;
	input_is_infinite_dffe21_wo <= input_is_infinite_dffe21;
	input_is_infinite_dffe22_wi <= input_is_infinite_dffe2_wo;
	input_is_infinite_dffe22_wo <= input_is_infinite_dffe22_wi;
	input_is_infinite_dffe23_wi <= input_is_infinite_dffe21_wo;
	input_is_infinite_dffe23_wo <= input_is_infinite_dffe23_wi;
	input_is_infinite_dffe25_wi <= input_is_infinite_dffe1_wo;
	input_is_infinite_dffe25_wo <= input_is_infinite_dffe25_wi;
	input_is_infinite_dffe26_wi <= input_is_infinite_dffe23_wo;
	input_is_infinite_dffe26_wo <= input_is_infinite_dffe26_wi;
	input_is_infinite_dffe27_wi <= input_is_infinite_dffe22_wo;
	input_is_infinite_dffe27_wo <= input_is_infinite_dffe27_wi;
	input_is_infinite_dffe2_wi <= input_is_infinite_dffe25_wo;
	input_is_infinite_dffe2_wo <= input_is_infinite_dffe2;
	input_is_infinite_dffe31_wi <= input_is_infinite_dffe26_wo;
	input_is_infinite_dffe31_wo <= input_is_infinite_dffe31;
	input_is_infinite_dffe32_wi <= input_is_infinite_dffe31_wo;
	input_is_infinite_dffe32_wo <= input_is_infinite_dffe32_wi;
	input_is_infinite_dffe33_wi <= input_is_infinite_dffe32_wo;
	input_is_infinite_dffe33_wo <= input_is_infinite_dffe33_wi;
	input_is_infinite_dffe3_wi <= input_is_infinite_dffe33_wo;
	input_is_infinite_dffe3_wo <= input_is_infinite_dffe3;
	input_is_infinite_dffe41_wi <= input_is_infinite_dffe42_wo;
	input_is_infinite_dffe41_wo <= input_is_infinite_dffe41_wi;
	input_is_infinite_dffe42_wi <= input_is_infinite_dffe3_wo;
	input_is_infinite_dffe42_wo <= input_is_infinite_dffe42_wi;
	input_is_infinite_dffe4_wi <= input_is_infinite_dffe41_wo;
	input_is_infinite_dffe4_wo <= input_is_infinite_dffe4;
	input_is_nan_dffe13_wi <= (input_dataa_nan_dffe12_wo OR input_datab_nan_dffe12_wo);
	input_is_nan_dffe13_wo <= input_is_nan_dffe13_wi;
	input_is_nan_dffe14_wi <= input_is_nan_dffe13_wo;
	input_is_nan_dffe14_wo <= input_is_nan_dffe14_wi;
	input_is_nan_dffe15_wi <= input_is_nan_dffe14_wo;
	input_is_nan_dffe15_wo <= input_is_nan_dffe15_wi;
	input_is_nan_dffe1_wi <= input_is_nan_dffe15_wo;
	input_is_nan_dffe1_wo <= input_is_nan_dffe1;
	input_is_nan_dffe21_wi <= input_is_nan_dffe27_wo;
	input_is_nan_dffe21_wo <= input_is_nan_dffe21;
	input_is_nan_dffe22_wi <= input_is_nan_dffe2_wo;
	input_is_nan_dffe22_wo <= input_is_nan_dffe22_wi;
	input_is_nan_dffe23_wi <= input_is_nan_dffe21_wo;
	input_is_nan_dffe23_wo <= input_is_nan_dffe23_wi;
	input_is_nan_dffe25_wi <= input_is_nan_dffe1_wo;
	input_is_nan_dffe25_wo <= input_is_nan_dffe25_wi;
	input_is_nan_dffe26_wi <= input_is_nan_dffe23_wo;
	input_is_nan_dffe26_wo <= input_is_nan_dffe26_wi;
	input_is_nan_dffe27_wi <= input_is_nan_dffe22_wo;
	input_is_nan_dffe27_wo <= input_is_nan_dffe27_wi;
	input_is_nan_dffe2_wi <= input_is_nan_dffe25_wo;
	input_is_nan_dffe2_wo <= input_is_nan_dffe2;
	input_is_nan_dffe31_wi <= input_is_nan_dffe26_wo;
	input_is_nan_dffe31_wo <= input_is_nan_dffe31;
	input_is_nan_dffe32_wi <= input_is_nan_dffe31_wo;
	input_is_nan_dffe32_wo <= input_is_nan_dffe32_wi;
	input_is_nan_dffe33_wi <= input_is_nan_dffe32_wo;
	input_is_nan_dffe33_wo <= input_is_nan_dffe33_wi;
	input_is_nan_dffe3_wi <= input_is_nan_dffe33_wo;
	input_is_nan_dffe3_wo <= input_is_nan_dffe3;
	input_is_nan_dffe41_wi <= input_is_nan_dffe42_wo;
	input_is_nan_dffe41_wo <= input_is_nan_dffe41_wi;
	input_is_nan_dffe42_wi <= input_is_nan_dffe3_wo;
	input_is_nan_dffe42_wo <= input_is_nan_dffe42_wi;
	input_is_nan_dffe4_wi <= input_is_nan_dffe41_wo;
	input_is_nan_dffe4_wo <= input_is_nan_dffe4;
	man_2comp_res_dataa_w <= ( pos_sign_bit_ext & datab_man_dffe1_wo);
	man_2comp_res_datab_w <= ( pos_sign_bit_ext & dataa_man_dffe1_wo);
	man_2comp_res_w <= ( wire_man_2comp_res_lower_w_lg_w_lg_w_lg_cout381w382w383w & wire_man_2comp_res_lower_result);
	man_a_not_zero_w <= ( wire_w_lg_w_dataa_range213w214w & wire_w_lg_w_dataa_range207w208w & wire_w_lg_w_dataa_range201w202w & wire_w_lg_w_dataa_range195w196w & wire_w_lg_w_dataa_range189w190w & wire_w_lg_w_dataa_range183w184w & wire_w_lg_w_dataa_range177w178w & wire_w_lg_w_dataa_range171w172w & wire_w_lg_w_dataa_range165w166w & wire_w_lg_w_dataa_range159w160w & wire_w_lg_w_dataa_range153w154w & wire_w_lg_w_dataa_range147w148w & wire_w_lg_w_dataa_range141w142w & wire_w_lg_w_dataa_range135w136w & wire_w_lg_w_dataa_range129w130w & wire_w_lg_w_dataa_range123w124w & wire_w_lg_w_dataa_range117w118w & wire_w_lg_w_dataa_range111w112w & wire_w_lg_w_dataa_range105w106w & wire_w_lg_w_dataa_range99w100w & wire_w_lg_w_dataa_range93w94w & wire_w_lg_w_dataa_range87w88w & dataa(0));
	man_add_sub_dataa_w <= ( pos_sign_bit_ext & dataa_man_dffe1_wo);
	man_add_sub_datab_w <= ( pos_sign_bit_ext & datab_man_dffe1_wo);
	man_add_sub_res_mag_dffe21_wi <= man_res_mag_w2;
	man_add_sub_res_mag_dffe21_wo <= man_add_sub_res_mag_dffe21;
	man_add_sub_res_mag_dffe23_wi <= man_add_sub_res_mag_dffe21_wo;
	man_add_sub_res_mag_dffe23_wo <= man_add_sub_res_mag_dffe23_wi;
	man_add_sub_res_mag_dffe26_wi <= man_add_sub_res_mag_dffe23_wo;
	man_add_sub_res_mag_dffe26_wo <= man_add_sub_res_mag_dffe26_wi;
	man_add_sub_res_mag_dffe27_wi <= man_add_sub_res_mag_w2;
	man_add_sub_res_mag_dffe27_wo <= man_add_sub_res_mag_dffe27_wi;
	man_add_sub_res_mag_w2 <= (wire_w_lg_w_man_add_sub_w_range386w393w OR wire_w_lg_w_lg_w_man_add_sub_w_range386w389w392w);
	man_add_sub_res_sign_dffe21_wo <= man_add_sub_res_sign_dffe21;
	man_add_sub_res_sign_dffe23_wi <= man_add_sub_res_sign_dffe21_wo;
	man_add_sub_res_sign_dffe23_wo <= man_add_sub_res_sign_dffe23_wi;
	man_add_sub_res_sign_dffe26_wi <= man_add_sub_res_sign_dffe23_wo;
	man_add_sub_res_sign_dffe26_wo <= man_add_sub_res_sign_dffe26_wi;
	man_add_sub_res_sign_dffe27_wi <= man_add_sub_res_sign_w2;
	man_add_sub_res_sign_dffe27_wo <= man_add_sub_res_sign_dffe27_wi;
	man_add_sub_res_sign_w2 <= (wire_w_lg_need_complement_dffe22_wo390w(0) OR (wire_w_lg_need_complement_dffe22_wo387w(0) AND man_add_sub_w(27)));
	man_add_sub_w <= ( wire_man_add_sub_lower_w_lg_w_lg_w_lg_cout368w369w370w & wire_man_add_sub_lower_result);
	man_all_zeros_w <= (OTHERS => '0');
	man_b_not_zero_w <= ( wire_w_lg_w_datab_range216w217w & wire_w_lg_w_datab_range210w211w & wire_w_lg_w_datab_range204w205w & wire_w_lg_w_datab_range198w199w & wire_w_lg_w_datab_range192w193w & wire_w_lg_w_datab_range186w187w & wire_w_lg_w_datab_range180w181w & wire_w_lg_w_datab_range174w175w & wire_w_lg_w_datab_range168w169w & wire_w_lg_w_datab_range162w163w & wire_w_lg_w_datab_range156w157w & wire_w_lg_w_datab_range150w151w & wire_w_lg_w_datab_range144w145w & wire_w_lg_w_datab_range138w139w & wire_w_lg_w_datab_range132w133w & wire_w_lg_w_datab_range126w127w & wire_w_lg_w_datab_range120w121w & wire_w_lg_w_datab_range114w115w & wire_w_lg_w_datab_range108w109w & wire_w_lg_w_datab_range102w103w & wire_w_lg_w_datab_range96w97w & wire_w_lg_w_datab_range90w91w & datab(0));
	man_dffe31_wo <= man_dffe31;
	man_intermediate_res_w <= ( "00" & man_res_w3);
	man_leading_zeros_cnt_w <= man_leading_zeros_dffe31_wo;
	man_leading_zeros_dffe31_wi <= (NOT wire_leading_zeroes_cnt_q);
	man_leading_zeros_dffe31_wo <= man_leading_zeros_dffe31;
	man_nan_w <= "10000000000000000000000";
	man_out_dffe5_wi <= (wire_w_lg_force_nan_w666w OR wire_w_lg_w_lg_force_nan_w644w665w);
	man_out_dffe5_wo <= man_out_dffe5;
	man_res_dffe4_wi <= man_rounded_res_w;
	man_res_dffe4_wo <= man_res_dffe4;
	man_res_is_not_zero_dffe31_wi <= man_res_not_zero_dffe26_wo;
	man_res_is_not_zero_dffe31_wo <= man_res_is_not_zero_dffe31;
	man_res_is_not_zero_dffe32_wi <= man_res_is_not_zero_dffe31_wo;
	man_res_is_not_zero_dffe32_wo <= man_res_is_not_zero_dffe32_wi;
	man_res_is_not_zero_dffe33_wi <= man_res_is_not_zero_dffe32_wo;
	man_res_is_not_zero_dffe33_wo <= man_res_is_not_zero_dffe33_wi;
	man_res_is_not_zero_dffe3_wi <= man_res_is_not_zero_dffe33_wo;
	man_res_is_not_zero_dffe3_wo <= man_res_is_not_zero_dffe3;
	man_res_is_not_zero_dffe41_wi <= man_res_is_not_zero_dffe42_wo;
	man_res_is_not_zero_dffe41_wo <= man_res_is_not_zero_dffe41_wi;
	man_res_is_not_zero_dffe42_wi <= man_res_is_not_zero_dffe3_wo;
	man_res_is_not_zero_dffe42_wo <= man_res_is_not_zero_dffe42_wi;
	man_res_is_not_zero_dffe4_wi <= man_res_is_not_zero_dffe41_wo;
	man_res_is_not_zero_dffe4_wo <= man_res_is_not_zero_dffe4;
	man_res_mag_w2 <= (wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w428w OR wire_w426w);
	man_res_not_zero_dffe23_wi <= man_res_not_zero_w2(24);
	man_res_not_zero_dffe23_wo <= man_res_not_zero_dffe23_wi;
	man_res_not_zero_dffe26_wi <= man_res_not_zero_dffe23_wo;
	man_res_not_zero_dffe26_wo <= man_res_not_zero_dffe26_wi;
	man_res_not_zero_w2 <= ( wire_w_lg_w_man_res_not_zero_w2_range501w503w & wire_w_lg_w_man_res_not_zero_w2_range498w500w & wire_w_lg_w_man_res_not_zero_w2_range495w497w & wire_w_lg_w_man_res_not_zero_w2_range492w494w & wire_w_lg_w_man_res_not_zero_w2_range489w491w & wire_w_lg_w_man_res_not_zero_w2_range486w488w & wire_w_lg_w_man_res_not_zero_w2_range483w485w & wire_w_lg_w_man_res_not_zero_w2_range480w482w & wire_w_lg_w_man_res_not_zero_w2_range477w479w & wire_w_lg_w_man_res_not_zero_w2_range474w476w & wire_w_lg_w_man_res_not_zero_w2_range471w473w & wire_w_lg_w_man_res_not_zero_w2_range468w470w & wire_w_lg_w_man_res_not_zero_w2_range465w467w & wire_w_lg_w_man_res_not_zero_w2_range462w464w & wire_w_lg_w_man_res_not_zero_w2_range459w461w & wire_w_lg_w_man_res_not_zero_w2_range456w458w & wire_w_lg_w_man_res_not_zero_w2_range453w455w & wire_w_lg_w_man_res_not_zero_w2_range450w452w & wire_w_lg_w_man_res_not_zero_w2_range447w449w & wire_w_lg_w_man_res_not_zero_w2_range444w446w & wire_w_lg_w_man_res_not_zero_w2_range441w443w & wire_w_lg_w_man_res_not_zero_w2_range438w440w & wire_w_lg_w_man_res_not_zero_w2_range435w437w & wire_w_lg_w_man_res_not_zero_w2_range431w434w & man_add_sub_res_mag_dffe21_wo(1));
	man_res_rounding_add_sub_datab_w <= ( "0000000000000000000000000" & man_rounding_add_value_w);
	man_res_rounding_add_sub_w <= ( wire_man_res_rounding_add_sub_lower_w_lg_w_lg_w_lg_cout594w595w596w & wire_man_res_rounding_add_sub_lower_result);
	man_res_w3 <= wire_lbarrel_shift_result(25 DOWNTO 2);
	man_rounded_res_w <= (wire_w_lg_w_man_res_rounding_add_sub_w_range599w603w OR wire_w601w);
	man_rounding_add_value_w <= (round_bit_dffe3_wo AND (sticky_bit_dffe3_wo OR guard_bit_dffe3_wo));
	man_smaller_dffe13_wi <= man_smaller_w;
	man_smaller_dffe13_wo <= man_smaller_dffe13_wi;
	man_smaller_w <= (wire_w_lg_exp_amb_mux_w279w OR wire_w_lg_w_lg_exp_amb_mux_w275w278w);
	need_complement_dffe22_wi <= need_complement_dffe2_wo;
	need_complement_dffe22_wo <= need_complement_dffe22_wi;
	need_complement_dffe2_wi <= dataa_sign_dffe25_wo;
	need_complement_dffe2_wo <= need_complement_dffe2;
	pos_sign_bit_ext <= (OTHERS => '0');
	priority_encoder_1pads_w <= (OTHERS => '1');
	result <= ( sign_out_dffe5_wo & exp_out_dffe5_wo & man_out_dffe5_wo);
	round_bit_dffe21_wi <= round_bit_w;
	round_bit_dffe21_wo <= round_bit_dffe21;
	round_bit_dffe23_wi <= round_bit_dffe21_wo;
	round_bit_dffe23_wo <= round_bit_dffe23_wi;
	round_bit_dffe26_wi <= round_bit_dffe23_wo;
	round_bit_dffe26_wo <= round_bit_dffe26_wi;
	round_bit_dffe31_wi <= round_bit_dffe26_wo;
	round_bit_dffe31_wo <= round_bit_dffe31;
	round_bit_dffe32_wi <= round_bit_dffe31_wo;
	round_bit_dffe32_wo <= round_bit_dffe32_wi;
	round_bit_dffe33_wi <= round_bit_dffe32_wo;
	round_bit_dffe33_wo <= round_bit_dffe33_wi;
	round_bit_dffe3_wi <= round_bit_dffe33_wo;
	round_bit_dffe3_wo <= round_bit_dffe3;
	round_bit_w <= ((((wire_w411w(0) AND man_add_sub_res_mag_dffe27_wo(0)) OR ((wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) AND man_add_sub_res_mag_dffe27_wo(25)) AND man_add_sub_res_mag_dffe27_wo(1))) OR (wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w405w(0) AND man_add_sub_res_mag_dffe27_wo(2))) OR ((man_add_sub_res_mag_dffe27_wo(26) AND man_add_sub_res_mag_dffe27_wo(25)) AND man_add_sub_res_mag_dffe27_wo(2)));
	rounded_res_infinity_dffe4_wi <= exp_rounded_res_infinity_w;
	rounded_res_infinity_dffe4_wo <= rounded_res_infinity_dffe4;
	rshift_distance_dffe13_wi <= rshift_distance_w;
	rshift_distance_dffe13_wo <= rshift_distance_dffe13_wi;
	rshift_distance_dffe14_wi <= rshift_distance_dffe13_wo;
	rshift_distance_dffe14_wo <= rshift_distance_dffe14_wi;
	rshift_distance_dffe15_wi <= rshift_distance_dffe14_wo;
	rshift_distance_dffe15_wo <= rshift_distance_dffe15_wi;
	rshift_distance_w <= (wire_w_lg_w_exp_diff_abs_exceed_max_w_range289w293w OR wire_w292w);
	sign_dffe31_wi <= ((man_res_not_zero_dffe26_wo AND man_add_sub_res_sign_dffe26_wo) OR wire_w_lg_w_lg_man_res_not_zero_dffe26_wo517w518w(0));
	sign_dffe31_wo <= sign_dffe31;
	sign_dffe32_wi <= sign_dffe31_wo;
	sign_dffe32_wo <= sign_dffe32_wi;
	sign_dffe33_wi <= sign_dffe32_wo;
	sign_dffe33_wo <= sign_dffe33_wi;
	sign_out_dffe5_wi <= (wire_w_lg_force_nan_w644w(0) AND ((force_infinity_w AND infinite_output_sign_dffe4_wo) OR wire_w_lg_w_lg_force_infinity_w643w668w(0)));
	sign_out_dffe5_wo <= sign_out_dffe5;
	sign_res_dffe3_wi <= sign_dffe33_wo;
	sign_res_dffe3_wo <= sign_res_dffe3;
	sign_res_dffe41_wi <= sign_res_dffe42_wo;
	sign_res_dffe41_wo <= sign_res_dffe41_wi;
	sign_res_dffe42_wi <= sign_res_dffe3_wo;
	sign_res_dffe42_wo <= sign_res_dffe42_wi;
	sign_res_dffe4_wi <= sign_res_dffe41_wo;
	sign_res_dffe4_wo <= sign_res_dffe4;
	sticky_bit_cnt_dataa_w <= ( "0" & rshift_distance_dffe15_wo);
	sticky_bit_cnt_datab_w <= ( "0" & wire_trailing_zeros_cnt_q);
	sticky_bit_cnt_res_w <= wire_add_sub3_result;
	sticky_bit_dffe1_wi <= wire_trailing_zeros_limit_comparator_agb;
	sticky_bit_dffe1_wo <= sticky_bit_dffe1;
	sticky_bit_dffe21_wi <= sticky_bit_w;
	sticky_bit_dffe21_wo <= sticky_bit_dffe21;
	sticky_bit_dffe22_wi <= sticky_bit_dffe2_wo;
	sticky_bit_dffe22_wo <= sticky_bit_dffe22_wi;
	sticky_bit_dffe23_wi <= sticky_bit_dffe21_wo;
	sticky_bit_dffe23_wo <= sticky_bit_dffe23_wi;
	sticky_bit_dffe25_wi <= sticky_bit_dffe1_wo;
	sticky_bit_dffe25_wo <= sticky_bit_dffe25_wi;
	sticky_bit_dffe26_wi <= sticky_bit_dffe23_wo;
	sticky_bit_dffe26_wo <= sticky_bit_dffe26_wi;
	sticky_bit_dffe27_wi <= sticky_bit_dffe22_wo;
	sticky_bit_dffe27_wo <= sticky_bit_dffe27_wi;
	sticky_bit_dffe2_wi <= sticky_bit_dffe25_wo;
	sticky_bit_dffe2_wo <= sticky_bit_dffe2;
	sticky_bit_dffe31_wi <= sticky_bit_dffe26_wo;
	sticky_bit_dffe31_wo <= sticky_bit_dffe31;
	sticky_bit_dffe32_wi <= sticky_bit_dffe31_wo;
	sticky_bit_dffe32_wo <= sticky_bit_dffe32_wi;
	sticky_bit_dffe33_wi <= sticky_bit_dffe32_wo;
	sticky_bit_dffe33_wo <= sticky_bit_dffe33_wi;
	sticky_bit_dffe3_wi <= sticky_bit_dffe33_wo;
	sticky_bit_dffe3_wo <= sticky_bit_dffe3;
	sticky_bit_w <= (((wire_w_lg_w411w421w(0) OR ((wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w396w(0) AND man_add_sub_res_mag_dffe27_wo(25)) AND wire_w_lg_sticky_bit_dffe27_wo416w(0))) OR (wire_w_lg_w_man_add_sub_res_mag_dffe27_wo_range395w405w(0) AND (wire_w_lg_sticky_bit_dffe27_wo416w(0) OR man_add_sub_res_mag_dffe27_wo(1)))) OR ((man_add_sub_res_mag_dffe27_wo(26) AND man_add_sub_res_mag_dffe27_wo(25)) AND (wire_w_lg_sticky_bit_dffe27_wo416w(0) OR man_add_sub_res_mag_dffe27_wo(1))));
	trailing_zeros_limit_w <= "000010";
	zero_man_sign_dffe21_wi <= zero_man_sign_dffe27_wo;
	zero_man_sign_dffe21_wo <= zero_man_sign_dffe21;
	zero_man_sign_dffe22_wi <= zero_man_sign_dffe2_wo;
	zero_man_sign_dffe22_wo <= zero_man_sign_dffe22_wi;
	zero_man_sign_dffe23_wi <= zero_man_sign_dffe21_wo;
	zero_man_sign_dffe23_wo <= zero_man_sign_dffe23_wi;
	zero_man_sign_dffe26_wi <= zero_man_sign_dffe23_wo;
	zero_man_sign_dffe26_wo <= zero_man_sign_dffe26_wi;
	zero_man_sign_dffe27_wi <= zero_man_sign_dffe22_wo;
	zero_man_sign_dffe27_wo <= zero_man_sign_dffe27_wi;
	zero_man_sign_dffe2_wi <= (dataa_sign_dffe25_wo AND add_sub_dffe25_wo);
	zero_man_sign_dffe2_wo <= zero_man_sign_dffe2;
	wire_w_aligned_dataa_exp_dffe15_wo_range315w <= aligned_dataa_exp_dffe15_wo(7 DOWNTO 0);
	wire_w_aligned_datab_exp_dffe15_wo_range313w <= aligned_datab_exp_dffe15_wo(7 DOWNTO 0);
	wire_w_dataa_range141w(0) <= dataa(10);
	wire_w_dataa_range147w(0) <= dataa(11);
	wire_w_dataa_range153w(0) <= dataa(12);
	wire_w_dataa_range159w(0) <= dataa(13);
	wire_w_dataa_range165w(0) <= dataa(14);
	wire_w_dataa_range171w(0) <= dataa(15);
	wire_w_dataa_range177w(0) <= dataa(16);
	wire_w_dataa_range183w(0) <= dataa(17);
	wire_w_dataa_range189w(0) <= dataa(18);
	wire_w_dataa_range195w(0) <= dataa(19);
	wire_w_dataa_range87w(0) <= dataa(1);
	wire_w_dataa_range201w(0) <= dataa(20);
	wire_w_dataa_range207w(0) <= dataa(21);
	wire_w_dataa_range213w(0) <= dataa(22);
	wire_w_dataa_range17w(0) <= dataa(24);
	wire_w_dataa_range27w(0) <= dataa(25);
	wire_w_dataa_range37w(0) <= dataa(26);
	wire_w_dataa_range47w(0) <= dataa(27);
	wire_w_dataa_range57w(0) <= dataa(28);
	wire_w_dataa_range67w(0) <= dataa(29);
	wire_w_dataa_range93w(0) <= dataa(2);
	wire_w_dataa_range77w(0) <= dataa(30);
	wire_w_dataa_range99w(0) <= dataa(3);
	wire_w_dataa_range105w(0) <= dataa(4);
	wire_w_dataa_range111w(0) <= dataa(5);
	wire_w_dataa_range117w(0) <= dataa(6);
	wire_w_dataa_range123w(0) <= dataa(7);
	wire_w_dataa_range129w(0) <= dataa(8);
	wire_w_dataa_range135w(0) <= dataa(9);
	wire_w_dataa_dffe11_wo_range242w <= dataa_dffe11_wo(22 DOWNTO 0);
	wire_w_dataa_dffe11_wo_range232w <= dataa_dffe11_wo(30 DOWNTO 23);
	wire_w_datab_range144w(0) <= datab(10);
	wire_w_datab_range150w(0) <= datab(11);
	wire_w_datab_range156w(0) <= datab(12);
	wire_w_datab_range162w(0) <= datab(13);
	wire_w_datab_range168w(0) <= datab(14);
	wire_w_datab_range174w(0) <= datab(15);
	wire_w_datab_range180w(0) <= datab(16);
	wire_w_datab_range186w(0) <= datab(17);
	wire_w_datab_range192w(0) <= datab(18);
	wire_w_datab_range198w(0) <= datab(19);
	wire_w_datab_range90w(0) <= datab(1);
	wire_w_datab_range204w(0) <= datab(20);
	wire_w_datab_range210w(0) <= datab(21);
	wire_w_datab_range216w(0) <= datab(22);
	wire_w_datab_range20w(0) <= datab(24);
	wire_w_datab_range30w(0) <= datab(25);
	wire_w_datab_range40w(0) <= datab(26);
	wire_w_datab_range50w(0) <= datab(27);
	wire_w_datab_range60w(0) <= datab(28);
	wire_w_datab_range70w(0) <= datab(29);
	wire_w_datab_range96w(0) <= datab(2);
	wire_w_datab_range80w(0) <= datab(30);
	wire_w_datab_range102w(0) <= datab(3);
	wire_w_datab_range108w(0) <= datab(4);
	wire_w_datab_range114w(0) <= datab(5);
	wire_w_datab_range120w(0) <= datab(6);
	wire_w_datab_range126w(0) <= datab(7);
	wire_w_datab_range132w(0) <= datab(8);
	wire_w_datab_range138w(0) <= datab(9);
	wire_w_datab_dffe11_wo_range261w <= datab_dffe11_wo(22 DOWNTO 0);
	wire_w_datab_dffe11_wo_range251w <= datab_dffe11_wo(30 DOWNTO 23);
	wire_w_exp_a_all_one_w_range7w(0) <= exp_a_all_one_w(0);
	wire_w_exp_a_all_one_w_range24w(0) <= exp_a_all_one_w(1);
	wire_w_exp_a_all_one_w_range34w(0) <= exp_a_all_one_w(2);
	wire_w_exp_a_all_one_w_range44w(0) <= exp_a_all_one_w(3);
	wire_w_exp_a_all_one_w_range54w(0) <= exp_a_all_one_w(4);
	wire_w_exp_a_all_one_w_range64w(0) <= exp_a_all_one_w(5);
	wire_w_exp_a_all_one_w_range74w(0) <= exp_a_all_one_w(6);
	wire_w_exp_a_all_one_w_range84w(0) <= exp_a_all_one_w(7);
	wire_w_exp_a_not_zero_w_range2w(0) <= exp_a_not_zero_w(0);
	wire_w_exp_a_not_zero_w_range19w(0) <= exp_a_not_zero_w(1);
	wire_w_exp_a_not_zero_w_range29w(0) <= exp_a_not_zero_w(2);
	wire_w_exp_a_not_zero_w_range39w(0) <= exp_a_not_zero_w(3);
	wire_w_exp_a_not_zero_w_range49w(0) <= exp_a_not_zero_w(4);
	wire_w_exp_a_not_zero_w_range59w(0) <= exp_a_not_zero_w(5);
	wire_w_exp_a_not_zero_w_range69w(0) <= exp_a_not_zero_w(6);
	wire_w_exp_adjustment2_add_sub_w_range532w(0) <= exp_adjustment2_add_sub_w(1);
	wire_w_exp_adjustment2_add_sub_w_range535w(0) <= exp_adjustment2_add_sub_w(2);
	wire_w_exp_adjustment2_add_sub_w_range538w(0) <= exp_adjustment2_add_sub_w(3);
	wire_w_exp_adjustment2_add_sub_w_range541w(0) <= exp_adjustment2_add_sub_w(4);
	wire_w_exp_adjustment2_add_sub_w_range544w(0) <= exp_adjustment2_add_sub_w(5);
	wire_w_exp_adjustment2_add_sub_w_range547w(0) <= exp_adjustment2_add_sub_w(6);
	wire_w_exp_adjustment2_add_sub_w_range571w <= exp_adjustment2_add_sub_w(7 DOWNTO 0);
	wire_w_exp_adjustment2_add_sub_w_range550w(0) <= exp_adjustment2_add_sub_w(7);
	wire_w_exp_adjustment2_add_sub_w_range525w(0) <= exp_adjustment2_add_sub_w(8);
	wire_w_exp_amb_w_range274w <= exp_amb_w(7 DOWNTO 0);
	wire_w_exp_b_all_one_w_range9w(0) <= exp_b_all_one_w(0);
	wire_w_exp_b_all_one_w_range26w(0) <= exp_b_all_one_w(1);
	wire_w_exp_b_all_one_w_range36w(0) <= exp_b_all_one_w(2);
	wire_w_exp_b_all_one_w_range46w(0) <= exp_b_all_one_w(3);
	wire_w_exp_b_all_one_w_range56w(0) <= exp_b_all_one_w(4);
	wire_w_exp_b_all_one_w_range66w(0) <= exp_b_all_one_w(5);
	wire_w_exp_b_all_one_w_range76w(0) <= exp_b_all_one_w(6);
	wire_w_exp_b_all_one_w_range86w(0) <= exp_b_all_one_w(7);
	wire_w_exp_b_not_zero_w_range5w(0) <= exp_b_not_zero_w(0);
	wire_w_exp_b_not_zero_w_range22w(0) <= exp_b_not_zero_w(1);
	wire_w_exp_b_not_zero_w_range32w(0) <= exp_b_not_zero_w(2);
	wire_w_exp_b_not_zero_w_range42w(0) <= exp_b_not_zero_w(3);
	wire_w_exp_b_not_zero_w_range52w(0) <= exp_b_not_zero_w(4);
	wire_w_exp_b_not_zero_w_range62w(0) <= exp_b_not_zero_w(5);
	wire_w_exp_b_not_zero_w_range72w(0) <= exp_b_not_zero_w(6);
	wire_w_exp_bma_w_range272w <= exp_bma_w(7 DOWNTO 0);
	wire_w_exp_diff_abs_exceed_max_w_range282w(0) <= exp_diff_abs_exceed_max_w(0);
	wire_w_exp_diff_abs_exceed_max_w_range286w(0) <= exp_diff_abs_exceed_max_w(1);
	wire_w_exp_diff_abs_exceed_max_w_range289w(0) <= exp_diff_abs_exceed_max_w(2);
	wire_w_exp_diff_abs_w_range290w <= exp_diff_abs_w(4 DOWNTO 0);
	wire_w_exp_diff_abs_w_range284w(0) <= exp_diff_abs_w(6);
	wire_w_exp_diff_abs_w_range287w(0) <= exp_diff_abs_w(7);
	wire_w_exp_res_max_w_range554w(0) <= exp_res_max_w(0);
	wire_w_exp_res_max_w_range557w(0) <= exp_res_max_w(1);
	wire_w_exp_res_max_w_range559w(0) <= exp_res_max_w(2);
	wire_w_exp_res_max_w_range561w(0) <= exp_res_max_w(3);
	wire_w_exp_res_max_w_range563w(0) <= exp_res_max_w(4);
	wire_w_exp_res_max_w_range565w(0) <= exp_res_max_w(5);
	wire_w_exp_res_max_w_range567w(0) <= exp_res_max_w(6);
	wire_w_exp_res_max_w_range569w(0) <= exp_res_max_w(7);
	wire_w_exp_res_not_zero_w_range530w(0) <= exp_res_not_zero_w(0);
	wire_w_exp_res_not_zero_w_range534w(0) <= exp_res_not_zero_w(1);
	wire_w_exp_res_not_zero_w_range537w(0) <= exp_res_not_zero_w(2);
	wire_w_exp_res_not_zero_w_range540w(0) <= exp_res_not_zero_w(3);
	wire_w_exp_res_not_zero_w_range543w(0) <= exp_res_not_zero_w(4);
	wire_w_exp_res_not_zero_w_range546w(0) <= exp_res_not_zero_w(5);
	wire_w_exp_res_not_zero_w_range549w(0) <= exp_res_not_zero_w(6);
	wire_w_exp_res_not_zero_w_range552w(0) <= exp_res_not_zero_w(7);
	wire_w_exp_rounded_res_max_w_range615w(0) <= exp_rounded_res_max_w(0);
	wire_w_exp_rounded_res_max_w_range619w(0) <= exp_rounded_res_max_w(1);
	wire_w_exp_rounded_res_max_w_range622w(0) <= exp_rounded_res_max_w(2);
	wire_w_exp_rounded_res_max_w_range625w(0) <= exp_rounded_res_max_w(3);
	wire_w_exp_rounded_res_max_w_range628w(0) <= exp_rounded_res_max_w(4);
	wire_w_exp_rounded_res_max_w_range631w(0) <= exp_rounded_res_max_w(5);
	wire_w_exp_rounded_res_max_w_range634w(0) <= exp_rounded_res_max_w(6);
	wire_w_exp_rounded_res_w_range617w(0) <= exp_rounded_res_w(1);
	wire_w_exp_rounded_res_w_range620w(0) <= exp_rounded_res_w(2);
	wire_w_exp_rounded_res_w_range623w(0) <= exp_rounded_res_w(3);
	wire_w_exp_rounded_res_w_range626w(0) <= exp_rounded_res_w(4);
	wire_w_exp_rounded_res_w_range629w(0) <= exp_rounded_res_w(5);
	wire_w_exp_rounded_res_w_range632w(0) <= exp_rounded_res_w(6);
	wire_w_exp_rounded_res_w_range635w(0) <= exp_rounded_res_w(7);
	wire_w_man_a_not_zero_w_range12w(0) <= man_a_not_zero_w(0);
	wire_w_man_a_not_zero_w_range143w(0) <= man_a_not_zero_w(10);
	wire_w_man_a_not_zero_w_range149w(0) <= man_a_not_zero_w(11);
	wire_w_man_a_not_zero_w_range155w(0) <= man_a_not_zero_w(12);
	wire_w_man_a_not_zero_w_range161w(0) <= man_a_not_zero_w(13);
	wire_w_man_a_not_zero_w_range167w(0) <= man_a_not_zero_w(14);
	wire_w_man_a_not_zero_w_range173w(0) <= man_a_not_zero_w(15);
	wire_w_man_a_not_zero_w_range179w(0) <= man_a_not_zero_w(16);
	wire_w_man_a_not_zero_w_range185w(0) <= man_a_not_zero_w(17);
	wire_w_man_a_not_zero_w_range191w(0) <= man_a_not_zero_w(18);
	wire_w_man_a_not_zero_w_range197w(0) <= man_a_not_zero_w(19);
	wire_w_man_a_not_zero_w_range89w(0) <= man_a_not_zero_w(1);
	wire_w_man_a_not_zero_w_range203w(0) <= man_a_not_zero_w(20);
	wire_w_man_a_not_zero_w_range209w(0) <= man_a_not_zero_w(21);
	wire_w_man_a_not_zero_w_range215w(0) <= man_a_not_zero_w(22);
	wire_w_man_a_not_zero_w_range95w(0) <= man_a_not_zero_w(2);
	wire_w_man_a_not_zero_w_range101w(0) <= man_a_not_zero_w(3);
	wire_w_man_a_not_zero_w_range107w(0) <= man_a_not_zero_w(4);
	wire_w_man_a_not_zero_w_range113w(0) <= man_a_not_zero_w(5);
	wire_w_man_a_not_zero_w_range119w(0) <= man_a_not_zero_w(6);
	wire_w_man_a_not_zero_w_range125w(0) <= man_a_not_zero_w(7);
	wire_w_man_a_not_zero_w_range131w(0) <= man_a_not_zero_w(8);
	wire_w_man_a_not_zero_w_range137w(0) <= man_a_not_zero_w(9);
	wire_w_man_add_sub_res_mag_dffe21_wo_range457w(0) <= man_add_sub_res_mag_dffe21_wo(10);
	wire_w_man_add_sub_res_mag_dffe21_wo_range460w(0) <= man_add_sub_res_mag_dffe21_wo(11);
	wire_w_man_add_sub_res_mag_dffe21_wo_range463w(0) <= man_add_sub_res_mag_dffe21_wo(12);
	wire_w_man_add_sub_res_mag_dffe21_wo_range466w(0) <= man_add_sub_res_mag_dffe21_wo(13);
	wire_w_man_add_sub_res_mag_dffe21_wo_range469w(0) <= man_add_sub_res_mag_dffe21_wo(14);
	wire_w_man_add_sub_res_mag_dffe21_wo_range472w(0) <= man_add_sub_res_mag_dffe21_wo(15);
	wire_w_man_add_sub_res_mag_dffe21_wo_range475w(0) <= man_add_sub_res_mag_dffe21_wo(16);
	wire_w_man_add_sub_res_mag_dffe21_wo_range478w(0) <= man_add_sub_res_mag_dffe21_wo(17);
	wire_w_man_add_sub_res_mag_dffe21_wo_range481w(0) <= man_add_sub_res_mag_dffe21_wo(18);
	wire_w_man_add_sub_res_mag_dffe21_wo_range484w(0) <= man_add_sub_res_mag_dffe21_wo(19);
	wire_w_man_add_sub_res_mag_dffe21_wo_range487w(0) <= man_add_sub_res_mag_dffe21_wo(20);
	wire_w_man_add_sub_res_mag_dffe21_wo_range490w(0) <= man_add_sub_res_mag_dffe21_wo(21);
	wire_w_man_add_sub_res_mag_dffe21_wo_range493w(0) <= man_add_sub_res_mag_dffe21_wo(22);
	wire_w_man_add_sub_res_mag_dffe21_wo_range496w(0) <= man_add_sub_res_mag_dffe21_wo(23);
	wire_w_man_add_sub_res_mag_dffe21_wo_range499w(0) <= man_add_sub_res_mag_dffe21_wo(24);
	wire_w_man_add_sub_res_mag_dffe21_wo_range502w(0) <= man_add_sub_res_mag_dffe21_wo(25);
	wire_w_man_add_sub_res_mag_dffe21_wo_range433w(0) <= man_add_sub_res_mag_dffe21_wo(2);
	wire_w_man_add_sub_res_mag_dffe21_wo_range436w(0) <= man_add_sub_res_mag_dffe21_wo(3);
	wire_w_man_add_sub_res_mag_dffe21_wo_range439w(0) <= man_add_sub_res_mag_dffe21_wo(4);
	wire_w_man_add_sub_res_mag_dffe21_wo_range442w(0) <= man_add_sub_res_mag_dffe21_wo(5);
	wire_w_man_add_sub_res_mag_dffe21_wo_range445w(0) <= man_add_sub_res_mag_dffe21_wo(6);
	wire_w_man_add_sub_res_mag_dffe21_wo_range448w(0) <= man_add_sub_res_mag_dffe21_wo(7);
	wire_w_man_add_sub_res_mag_dffe21_wo_range451w(0) <= man_add_sub_res_mag_dffe21_wo(8);
	wire_w_man_add_sub_res_mag_dffe21_wo_range454w(0) <= man_add_sub_res_mag_dffe21_wo(9);
	wire_w_man_add_sub_res_mag_dffe27_wo_range410w(0) <= man_add_sub_res_mag_dffe27_wo(0);
	wire_w_man_add_sub_res_mag_dffe27_wo_range425w <= man_add_sub_res_mag_dffe27_wo(25 DOWNTO 0);
	wire_w_man_add_sub_res_mag_dffe27_wo_range401w(0) <= man_add_sub_res_mag_dffe27_wo(25);
	wire_w_man_add_sub_res_mag_dffe27_wo_range427w <= man_add_sub_res_mag_dffe27_wo(26 DOWNTO 1);
	wire_w_man_add_sub_res_mag_dffe27_wo_range395w(0) <= man_add_sub_res_mag_dffe27_wo(26);
	wire_w_man_add_sub_w_range386w(0) <= man_add_sub_w(27);
	wire_w_man_b_not_zero_w_range15w(0) <= man_b_not_zero_w(0);
	wire_w_man_b_not_zero_w_range146w(0) <= man_b_not_zero_w(10);
	wire_w_man_b_not_zero_w_range152w(0) <= man_b_not_zero_w(11);
	wire_w_man_b_not_zero_w_range158w(0) <= man_b_not_zero_w(12);
	wire_w_man_b_not_zero_w_range164w(0) <= man_b_not_zero_w(13);
	wire_w_man_b_not_zero_w_range170w(0) <= man_b_not_zero_w(14);
	wire_w_man_b_not_zero_w_range176w(0) <= man_b_not_zero_w(15);
	wire_w_man_b_not_zero_w_range182w(0) <= man_b_not_zero_w(16);
	wire_w_man_b_not_zero_w_range188w(0) <= man_b_not_zero_w(17);
	wire_w_man_b_not_zero_w_range194w(0) <= man_b_not_zero_w(18);
	wire_w_man_b_not_zero_w_range200w(0) <= man_b_not_zero_w(19);
	wire_w_man_b_not_zero_w_range92w(0) <= man_b_not_zero_w(1);
	wire_w_man_b_not_zero_w_range206w(0) <= man_b_not_zero_w(20);
	wire_w_man_b_not_zero_w_range212w(0) <= man_b_not_zero_w(21);
	wire_w_man_b_not_zero_w_range218w(0) <= man_b_not_zero_w(22);
	wire_w_man_b_not_zero_w_range98w(0) <= man_b_not_zero_w(2);
	wire_w_man_b_not_zero_w_range104w(0) <= man_b_not_zero_w(3);
	wire_w_man_b_not_zero_w_range110w(0) <= man_b_not_zero_w(4);
	wire_w_man_b_not_zero_w_range116w(0) <= man_b_not_zero_w(5);
	wire_w_man_b_not_zero_w_range122w(0) <= man_b_not_zero_w(6);
	wire_w_man_b_not_zero_w_range128w(0) <= man_b_not_zero_w(7);
	wire_w_man_b_not_zero_w_range134w(0) <= man_b_not_zero_w(8);
	wire_w_man_b_not_zero_w_range140w(0) <= man_b_not_zero_w(9);
	wire_w_man_res_not_zero_w2_range431w(0) <= man_res_not_zero_w2(0);
	wire_w_man_res_not_zero_w2_range462w(0) <= man_res_not_zero_w2(10);
	wire_w_man_res_not_zero_w2_range465w(0) <= man_res_not_zero_w2(11);
	wire_w_man_res_not_zero_w2_range468w(0) <= man_res_not_zero_w2(12);
	wire_w_man_res_not_zero_w2_range471w(0) <= man_res_not_zero_w2(13);
	wire_w_man_res_not_zero_w2_range474w(0) <= man_res_not_zero_w2(14);
	wire_w_man_res_not_zero_w2_range477w(0) <= man_res_not_zero_w2(15);
	wire_w_man_res_not_zero_w2_range480w(0) <= man_res_not_zero_w2(16);
	wire_w_man_res_not_zero_w2_range483w(0) <= man_res_not_zero_w2(17);
	wire_w_man_res_not_zero_w2_range486w(0) <= man_res_not_zero_w2(18);
	wire_w_man_res_not_zero_w2_range489w(0) <= man_res_not_zero_w2(19);
	wire_w_man_res_not_zero_w2_range435w(0) <= man_res_not_zero_w2(1);
	wire_w_man_res_not_zero_w2_range492w(0) <= man_res_not_zero_w2(20);
	wire_w_man_res_not_zero_w2_range495w(0) <= man_res_not_zero_w2(21);
	wire_w_man_res_not_zero_w2_range498w(0) <= man_res_not_zero_w2(22);
	wire_w_man_res_not_zero_w2_range501w(0) <= man_res_not_zero_w2(23);
	wire_w_man_res_not_zero_w2_range438w(0) <= man_res_not_zero_w2(2);
	wire_w_man_res_not_zero_w2_range441w(0) <= man_res_not_zero_w2(3);
	wire_w_man_res_not_zero_w2_range444w(0) <= man_res_not_zero_w2(4);
	wire_w_man_res_not_zero_w2_range447w(0) <= man_res_not_zero_w2(5);
	wire_w_man_res_not_zero_w2_range450w(0) <= man_res_not_zero_w2(6);
	wire_w_man_res_not_zero_w2_range453w(0) <= man_res_not_zero_w2(7);
	wire_w_man_res_not_zero_w2_range456w(0) <= man_res_not_zero_w2(8);
	wire_w_man_res_not_zero_w2_range459w(0) <= man_res_not_zero_w2(9);
	wire_w_man_res_rounding_add_sub_w_range598w <= man_res_rounding_add_sub_w(22 DOWNTO 0);
	wire_w_man_res_rounding_add_sub_w_range602w <= man_res_rounding_add_sub_w(23 DOWNTO 1);
	wire_w_man_res_rounding_add_sub_w_range599w(0) <= man_res_rounding_add_sub_w(24);
	lbarrel_shift :  addSub_altbarrel_shift_35e
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => man_dffe31_wo,
		distance => man_leading_zeros_cnt_w,
		result => wire_lbarrel_shift_result
	  );
	wire_rbarrel_shift_data <= ( man_smaller_dffe13_wo & "00");
	rbarrel_shift :  addSub_altbarrel_shift_olb
	  PORT MAP ( 
		data => wire_rbarrel_shift_data,
		distance => rshift_distance_dffe13_wo,
		result => wire_rbarrel_shift_result
	  );
	wire_leading_zeroes_cnt_data <= ( man_add_sub_res_mag_dffe21_wo(25 DOWNTO 1) & "1" & "000000");
	leading_zeroes_cnt :  addSub_altpriority_encoder_qb6
	  PORT MAP ( 
		data => wire_leading_zeroes_cnt_data,
		q => wire_leading_zeroes_cnt_q
	  );
	wire_trailing_zeros_cnt_data <= ( "111111111" & man_smaller_dffe13_wo(22 DOWNTO 0));
	trailing_zeros_cnt :  addSub_altpriority_encoder_e48
	  PORT MAP ( 
		data => wire_trailing_zeros_cnt_data,
		q => wire_trailing_zeros_cnt_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_sub_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_sub_dffe1 <= add_sub_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN both_inputs_are_infinite_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN both_inputs_are_infinite_dffe1 <= both_inputs_are_infinite_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN data_exp_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN data_exp_dffe1 <= data_exp_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_man_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_man_dffe1 <= dataa_man_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_sign_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_sign_dffe1 <= dataa_sign_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_man_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_man_dffe1 <= datab_man_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_sign_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_sign_dffe1 <= datab_sign_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN denormal_res_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN denormal_res_dffe3 <= denormal_res_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN denormal_res_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN denormal_res_dffe4 <= denormal_res_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_adj_dffe21 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_adj_dffe21 <= exp_adj_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_out_dffe5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_out_dffe5 <= exp_out_dffe5_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_res_dffe2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_res_dffe2 <= exp_res_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_res_dffe21 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_res_dffe21 <= exp_res_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_res_dffe3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_res_dffe3 <= exp_res_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_res_dffe4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_res_dffe4 <= exp_res_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe1 <= infinite_output_sign_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe2 <= infinite_output_sign_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe21 <= infinite_output_sign_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe3 <= infinite_output_sign_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe31 <= infinite_output_sign_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_output_sign_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_output_sign_dffe4 <= infinite_output_sign_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_res_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_res_dffe3 <= infinite_res_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_res_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_res_dffe4 <= infinite_res_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_magnitude_sub_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_magnitude_sub_dffe2 <= infinity_magnitude_sub_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_magnitude_sub_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_magnitude_sub_dffe21 <= infinity_magnitude_sub_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_magnitude_sub_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_magnitude_sub_dffe3 <= infinity_magnitude_sub_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_magnitude_sub_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_magnitude_sub_dffe31 <= infinity_magnitude_sub_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_magnitude_sub_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_magnitude_sub_dffe4 <= infinity_magnitude_sub_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe1 <= input_is_infinite_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe2 <= input_is_infinite_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe21 <= input_is_infinite_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe3 <= input_is_infinite_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe31 <= input_is_infinite_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinite_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinite_dffe4 <= input_is_infinite_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe1 <= input_is_nan_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe2 <= input_is_nan_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe21 <= input_is_nan_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe3 <= input_is_nan_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe31 <= input_is_nan_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe4 <= input_is_nan_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_add_sub_res_mag_dffe21 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_add_sub_res_mag_dffe21 <= man_add_sub_res_mag_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_add_sub_res_sign_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_add_sub_res_sign_dffe21 <= man_add_sub_res_sign_dffe27_wo;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe31 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe31 <= man_add_sub_res_mag_dffe26_wo;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_leading_zeros_dffe31 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_leading_zeros_dffe31 <= man_leading_zeros_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_out_dffe5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_out_dffe5 <= man_out_dffe5_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_res_dffe4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_res_dffe4 <= man_res_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_res_is_not_zero_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_res_is_not_zero_dffe3 <= man_res_is_not_zero_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_res_is_not_zero_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_res_is_not_zero_dffe31 <= man_res_is_not_zero_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_res_is_not_zero_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_res_is_not_zero_dffe4 <= man_res_is_not_zero_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN need_complement_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN need_complement_dffe2 <= need_complement_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_bit_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_bit_dffe21 <= round_bit_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_bit_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_bit_dffe3 <= round_bit_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_bit_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_bit_dffe31 <= round_bit_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rounded_res_infinity_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN rounded_res_infinity_dffe4 <= rounded_res_infinity_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe31 <= sign_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_out_dffe5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_out_dffe5 <= sign_out_dffe5_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_res_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_res_dffe3 <= sign_res_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_res_dffe4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_res_dffe4 <= sign_res_dffe4_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_bit_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_bit_dffe1 <= sticky_bit_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_bit_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_bit_dffe2 <= sticky_bit_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_bit_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_bit_dffe21 <= sticky_bit_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_bit_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_bit_dffe3 <= sticky_bit_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_bit_dffe31 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_bit_dffe31 <= sticky_bit_dffe31_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_man_sign_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_man_sign_dffe2 <= zero_man_sign_dffe2_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_man_sign_dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_man_sign_dffe21 <= zero_man_sign_dffe21_wi;
			END IF;
		END IF;
	END PROCESS;
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => aligned_dataa_exp_w,
		datab => aligned_datab_exp_w,
		result => wire_add_sub1_result
	  );
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => aligned_datab_exp_w,
		datab => aligned_dataa_exp_w,
		result => wire_add_sub2_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => sticky_bit_cnt_dataa_w,
		datab => sticky_bit_cnt_datab_w,
		result => wire_add_sub3_result
	  );
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => exp_adjustment_add_sub_dataa_w,
		datab => exp_adjustment_add_sub_datab_w,
		result => wire_add_sub4_result
	  );
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_adjustment2_add_sub_dataa_w,
		datab => exp_adjustment2_add_sub_datab_w,
		result => wire_add_sub5_result
	  );
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => exp_res_rounding_adder_dataa_w,
		datab => exp_rounding_adjustment_w,
		result => wire_add_sub6_result
	  );
	loop121 : FOR i IN 0 TO 13 GENERATE 
		wire_man_2comp_res_lower_w_lg_w_lg_cout381w382w(i) <= wire_man_2comp_res_lower_w_lg_cout381w(0) AND wire_man_2comp_res_upper0_result(i);
	END GENERATE loop121;
	loop122 : FOR i IN 0 TO 13 GENERATE 
		wire_man_2comp_res_lower_w_lg_cout380w(i) <= wire_man_2comp_res_lower_cout AND wire_man_2comp_res_upper1_result(i);
	END GENERATE loop122;
	wire_man_2comp_res_lower_w_lg_cout381w(0) <= NOT wire_man_2comp_res_lower_cout;
	loop123 : FOR i IN 0 TO 13 GENERATE 
		wire_man_2comp_res_lower_w_lg_w_lg_w_lg_cout381w382w383w(i) <= wire_man_2comp_res_lower_w_lg_w_lg_cout381w382w(i) OR wire_man_2comp_res_lower_w_lg_cout380w(i);
	END GENERATE loop123;
	man_2comp_res_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => borrow_w,
		clken => clk_en,
		clock => clock,
		cout => wire_man_2comp_res_lower_cout,
		dataa => man_2comp_res_dataa_w(13 DOWNTO 0),
		datab => man_2comp_res_datab_w(13 DOWNTO 0),
		result => wire_man_2comp_res_lower_result
	  );
	man_2comp_res_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => wire_gnd,
		clken => clk_en,
		clock => clock,
		dataa => man_2comp_res_dataa_w(27 DOWNTO 14),
		datab => man_2comp_res_datab_w(27 DOWNTO 14),
		result => wire_man_2comp_res_upper0_result
	  );
	man_2comp_res_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => wire_vcc,
		clken => clk_en,
		clock => clock,
		dataa => man_2comp_res_dataa_w(27 DOWNTO 14),
		datab => man_2comp_res_datab_w(27 DOWNTO 14),
		result => wire_man_2comp_res_upper1_result
	  );
	loop124 : FOR i IN 0 TO 13 GENERATE 
		wire_man_add_sub_lower_w_lg_w_lg_cout368w369w(i) <= wire_man_add_sub_lower_w_lg_cout368w(0) AND wire_man_add_sub_upper0_result(i);
	END GENERATE loop124;
	loop125 : FOR i IN 0 TO 13 GENERATE 
		wire_man_add_sub_lower_w_lg_cout367w(i) <= wire_man_add_sub_lower_cout AND wire_man_add_sub_upper1_result(i);
	END GENERATE loop125;
	wire_man_add_sub_lower_w_lg_cout368w(0) <= NOT wire_man_add_sub_lower_cout;
	loop126 : FOR i IN 0 TO 13 GENERATE 
		wire_man_add_sub_lower_w_lg_w_lg_w_lg_cout368w369w370w(i) <= wire_man_add_sub_lower_w_lg_w_lg_cout368w369w(i) OR wire_man_add_sub_lower_w_lg_cout367w(i);
	END GENERATE loop126;
	man_add_sub_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => borrow_w,
		clken => clk_en,
		clock => clock,
		cout => wire_man_add_sub_lower_cout,
		dataa => man_add_sub_dataa_w(13 DOWNTO 0),
		datab => man_add_sub_datab_w(13 DOWNTO 0),
		result => wire_man_add_sub_lower_result
	  );
	man_add_sub_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => wire_gnd,
		clken => clk_en,
		clock => clock,
		dataa => man_add_sub_dataa_w(27 DOWNTO 14),
		datab => man_add_sub_datab_w(27 DOWNTO 14),
		result => wire_man_add_sub_upper0_result
	  );
	man_add_sub_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 14,
		lpm_hint => "USE_WYS=ON"
	  )
	  PORT MAP ( 
		aclr => aclr,
		add_sub => add_sub_w2,
		cin => wire_vcc,
		clken => clk_en,
		clock => clock,
		dataa => man_add_sub_dataa_w(27 DOWNTO 14),
		datab => man_add_sub_datab_w(27 DOWNTO 14),
		result => wire_man_add_sub_upper1_result
	  );
	loop127 : FOR i IN 0 TO 12 GENERATE 
		wire_man_res_rounding_add_sub_lower_w_lg_w_lg_cout594w595w(i) <= wire_man_res_rounding_add_sub_lower_w_lg_cout594w(0) AND adder_upper_w(i);
	END GENERATE loop127;
	loop128 : FOR i IN 0 TO 12 GENERATE 
		wire_man_res_rounding_add_sub_lower_w_lg_cout593w(i) <= wire_man_res_rounding_add_sub_lower_cout AND wire_man_res_rounding_add_sub_upper1_result(i);
	END GENERATE loop128;
	wire_man_res_rounding_add_sub_lower_w_lg_cout594w(0) <= NOT wire_man_res_rounding_add_sub_lower_cout;
	loop129 : FOR i IN 0 TO 12 GENERATE 
		wire_man_res_rounding_add_sub_lower_w_lg_w_lg_w_lg_cout594w595w596w(i) <= wire_man_res_rounding_add_sub_lower_w_lg_w_lg_cout594w595w(i) OR wire_man_res_rounding_add_sub_lower_w_lg_cout593w(i);
	END GENERATE loop129;
	man_res_rounding_add_sub_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		cout => wire_man_res_rounding_add_sub_lower_cout,
		dataa => man_intermediate_res_w(12 DOWNTO 0),
		datab => man_res_rounding_add_sub_datab_w(12 DOWNTO 0),
		result => wire_man_res_rounding_add_sub_lower_result
	  );
	man_res_rounding_add_sub_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		cin => wire_vcc,
		dataa => man_intermediate_res_w(25 DOWNTO 13),
		datab => man_res_rounding_add_sub_datab_w(25 DOWNTO 13),
		result => wire_man_res_rounding_add_sub_upper1_result
	  );
	trailing_zeros_limit_comparator :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		agb => wire_trailing_zeros_limit_comparator_agb,
		dataa => sticky_bit_cnt_res_w,
		datab => trailing_zeros_limit_w
	  );

 END RTL; --addSub_altfp_add_sub_kdk
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY addSub IS
	PORT
	(
		add_sub		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END addSub;


ARCHITECTURE RTL OF addsub IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT addSub_altfp_add_sub_kdk
	PORT (
			add_sub	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	addSub_altfp_add_sub_kdk_component : addSub_altfp_add_sub_kdk
	PORT MAP (
		add_sub => add_sub,
		clock => clock,
		datab => datab,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIDTH_DATA NUMERIC "32"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: DIRECTION STRING "VARIABLE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: OPTIMIZE STRING "SPEED"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "7"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: add_sub 0 0 0 0 INPUT NODEFVAL "add_sub"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @add_sub 0 0 0 0 add_sub 0 0 0 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL addSub.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL addSub.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL addSub.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL addSub.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL addSub_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
