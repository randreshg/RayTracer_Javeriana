-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: convert.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" OPERATION="INT2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=32 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=32 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_altfp_convert 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_altsyncram 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_abs 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_decode 2013:06:12:18:03:43:SJ cbx_lpm_divide 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_stratixiii 2013:06:12:18:03:43:SJ cbx_stratixv 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = reg 68 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altbarrel_shift_tvf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END convert_altbarrel_shift_tvf;

 ARCHITECTURE RTL OF convert_altbarrel_shift_tvf IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w98w99w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w94w95w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w119w120w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w115w116w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w141w142w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w137w138w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w163w164w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w159w160w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w182w183w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w178w179w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w90w91w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w111w112w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w133w134w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w155w156w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w174w175w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range82w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range104w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range125w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range149w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range168w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w119w120w121w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w141w142w143w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w163w164w165w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w182w183w184w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w101w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w122w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w144w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w166w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w185w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w114w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w117w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w136w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w139w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w158w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w161w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w177w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w180w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range92w93w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w96w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range145w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range167w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range80w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range103w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range123w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range173w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range132w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w98w99w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w98w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w96w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w94w95w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w94w(0) AND wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range92w93w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w119w120w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w119w(0) AND wire_altbarrel_shift5_w117w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w115w116w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w115w(0) AND wire_altbarrel_shift5_w114w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w141w142w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w141w(0) AND wire_altbarrel_shift5_w139w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w137w138w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w137w(0) AND wire_altbarrel_shift5_w136w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w163w164w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w163w(0) AND wire_altbarrel_shift5_w161w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w159w160w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w159w(0) AND wire_altbarrel_shift5_w158w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w182w183w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w182w(0) AND wire_altbarrel_shift5_w180w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w178w179w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w178w(0) AND wire_altbarrel_shift5_w177w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w90w91w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w90w(0) AND wire_altbarrel_shift5_w_sbit_w_range80w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w111w112w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w111w(0) AND wire_altbarrel_shift5_w_sbit_w_range103w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w133w134w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w133w(0) AND wire_altbarrel_shift5_w_sbit_w_range123w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w155w156w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w155w(0) AND wire_altbarrel_shift5_w_sbit_w_range145w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w174w175w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w174w(0) AND wire_altbarrel_shift5_w_sbit_w_range167w(i);
	END GENERATE loop14;
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w98w(0) <= wire_altbarrel_shift5_w_sel_w_range85w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range82w97w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w94w(0) <= wire_altbarrel_shift5_w_sel_w_range85w(0) AND wire_altbarrel_shift5_w_dir_w_range82w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w119w(0) <= wire_altbarrel_shift5_w_sel_w_range106w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range104w118w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w115w(0) <= wire_altbarrel_shift5_w_sel_w_range106w(0) AND wire_altbarrel_shift5_w_dir_w_range104w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w141w(0) <= wire_altbarrel_shift5_w_sel_w_range128w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range125w140w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w137w(0) <= wire_altbarrel_shift5_w_sel_w_range128w(0) AND wire_altbarrel_shift5_w_dir_w_range125w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w163w(0) <= wire_altbarrel_shift5_w_sel_w_range151w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range149w162w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w159w(0) <= wire_altbarrel_shift5_w_sel_w_range151w(0) AND wire_altbarrel_shift5_w_dir_w_range149w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w182w(0) <= wire_altbarrel_shift5_w_sel_w_range170w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range168w181w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w178w(0) <= wire_altbarrel_shift5_w_sel_w_range170w(0) AND wire_altbarrel_shift5_w_dir_w_range168w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range82w97w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range82w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range104w118w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range104w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range125w140w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range125w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range149w162w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range149w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range168w181w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range168w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w90w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range85w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w111w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range106w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w133w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range128w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w155w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range151w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w174w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range170w(0);
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w98w99w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w94w95w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w119w120w121w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w119w120w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w115w116w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w141w142w143w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w141w142w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w137w138w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w163w164w165w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w163w164w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w159w160w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w182w183w184w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w182w183w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w178w179w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w101w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w90w91w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w122w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w119w120w121w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w111w112w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w144w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w141w142w143w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w133w134w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w166w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w163w164w165w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w155w156w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w185w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w182w183w184w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w174w175w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(1) & dir_w(3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper2d & smux_w(127 DOWNTO 96) & sbit_piper1d & smux_w(63 DOWNTO 0) & data);
	sel_w <= ( sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift5_w185w & wire_altbarrel_shift5_w166w & wire_altbarrel_shift5_w144w & wire_altbarrel_shift5_w122w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w98w99w100w101w);
	wire_altbarrel_shift5_w114w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_altbarrel_shift5_w117w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift5_w136w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_altbarrel_shift5_w139w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift5_w158w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_altbarrel_shift5_w161w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift5_w177w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_altbarrel_shift5_w180w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range92w93w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w96w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift5_w_dir_w_range82w(0) <= dir_w(0);
	wire_altbarrel_shift5_w_dir_w_range104w(0) <= dir_w(1);
	wire_altbarrel_shift5_w_dir_w_range125w(0) <= dir_w(2);
	wire_altbarrel_shift5_w_dir_w_range149w(0) <= dir_w(3);
	wire_altbarrel_shift5_w_dir_w_range168w(0) <= dir_w(4);
	wire_altbarrel_shift5_w_sbit_w_range145w <= sbit_w(127 DOWNTO 96);
	wire_altbarrel_shift5_w_sbit_w_range167w <= sbit_w(159 DOWNTO 128);
	wire_altbarrel_shift5_w_sbit_w_range80w <= sbit_w(31 DOWNTO 0);
	wire_altbarrel_shift5_w_sbit_w_range103w <= sbit_w(63 DOWNTO 32);
	wire_altbarrel_shift5_w_sbit_w_range123w <= sbit_w(95 DOWNTO 64);
	wire_altbarrel_shift5_w_sel_w_range85w(0) <= sel_w(0);
	wire_altbarrel_shift5_w_sel_w_range106w(0) <= sel_w(1);
	wire_altbarrel_shift5_w_sel_w_range128w(0) <= sel_w(2);
	wire_altbarrel_shift5_w_sel_w_range151w(0) <= sel_w(3);
	wire_altbarrel_shift5_w_sel_w_range170w(0) <= sel_w(4);
	wire_altbarrel_shift5_w_smux_w_range173w <= smux_w(159 DOWNTO 128);
	wire_altbarrel_shift5_w_smux_w_range132w <= smux_w(95 DOWNTO 64);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(4) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift5_w_smux_w_range132w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift5_w_smux_w_range173w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --convert_altbarrel_shift_tvf


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END convert_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF convert_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --convert_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END convert_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF convert_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero221w & wire_altpriority_encoder16_w_lg_w_lg_zero223w224w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  convert_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	wire_altpriority_encoder16_w_lg_w_lg_zero221w222w(0) <= wire_altpriority_encoder16_w_lg_zero221w(0) AND wire_altpriority_encoder16_q(0);
	wire_altpriority_encoder16_w_lg_zero223w(0) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder16_w_lg_zero221w(0) <= NOT wire_altpriority_encoder16_zero;
	wire_altpriority_encoder16_w_lg_w_lg_zero223w224w(0) <= wire_altpriority_encoder16_w_lg_zero223w(0) OR wire_altpriority_encoder16_w_lg_w_lg_zero221w222w(0);
	altpriority_encoder16 :  convert_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --convert_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END convert_altpriority_encoder_be8;

 ARCHITECTURE RTL OF convert_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero211w212w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero213w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero213w214w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero211w & wire_altpriority_encoder14_w_lg_w_lg_zero213w214w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  convert_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop25 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero211w212w(i) <= wire_altpriority_encoder14_w_lg_zero211w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero213w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop26;
	wire_altpriority_encoder14_w_lg_zero211w(0) <= NOT wire_altpriority_encoder14_zero;
	loop27 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero213w214w(i) <= wire_altpriority_encoder14_w_lg_zero213w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero211w212w(i);
	END GENERATE loop27;
	altpriority_encoder14 :  convert_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --convert_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END convert_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF convert_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero201w202w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero203w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero203w204w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero201w & wire_altpriority_encoder12_w_lg_w_lg_zero203w204w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  convert_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	loop28 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero201w202w(i) <= wire_altpriority_encoder12_w_lg_zero201w(0) AND wire_altpriority_encoder12_q(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_zero203w(i) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(i);
	END GENERATE loop29;
	wire_altpriority_encoder12_w_lg_zero201w(0) <= NOT wire_altpriority_encoder12_zero;
	loop30 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero203w204w(i) <= wire_altpriority_encoder12_w_lg_zero203w(i) OR wire_altpriority_encoder12_w_lg_w_lg_zero201w202w(i);
	END GENERATE loop30;
	altpriority_encoder12 :  convert_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --convert_altpriority_encoder_rf8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END convert_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF convert_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --convert_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END convert_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF convert_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero255w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  convert_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero255w & wire_altpriority_encoder22_w_lg_w_lg_zero257w258w);
	altpriority_encoder21 :  convert_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder21_q
	  );
	wire_altpriority_encoder22_w_lg_w_lg_zero255w256w(0) <= wire_altpriority_encoder22_w_lg_zero255w(0) AND wire_altpriority_encoder22_q(0);
	wire_altpriority_encoder22_w_lg_zero257w(0) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(0);
	wire_altpriority_encoder22_w_lg_zero255w(0) <= NOT wire_altpriority_encoder22_zero;
	wire_altpriority_encoder22_w_lg_w_lg_zero257w258w(0) <= wire_altpriority_encoder22_w_lg_zero257w(0) OR wire_altpriority_encoder22_w_lg_w_lg_zero255w256w(0);
	altpriority_encoder22 :  convert_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --convert_altpriority_encoder_6v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END convert_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF convert_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero246w247w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero248w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero248w249w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  convert_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero246w & wire_altpriority_encoder20_w_lg_w_lg_zero248w249w);
	altpriority_encoder19 :  convert_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop31 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero246w247w(i) <= wire_altpriority_encoder20_w_lg_zero246w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_zero248w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop32;
	wire_altpriority_encoder20_w_lg_zero246w(0) <= NOT wire_altpriority_encoder20_zero;
	loop33 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero248w249w(i) <= wire_altpriority_encoder20_w_lg_zero248w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero246w247w(i);
	END GENERATE loop33;
	altpriority_encoder20 :  convert_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --convert_altpriority_encoder_bv7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END convert_altpriority_encoder_r08;

 ARCHITECTURE RTL OF convert_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero237w238w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero239w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero239w240w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  convert_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  convert_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero237w & wire_altpriority_encoder18_w_lg_w_lg_zero239w240w);
	altpriority_encoder17 :  convert_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero237w238w(i) <= wire_altpriority_encoder18_w_lg_zero237w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_zero239w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop35;
	wire_altpriority_encoder18_w_lg_zero237w(0) <= NOT wire_altpriority_encoder18_zero;
	loop36 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero239w240w(i) <= wire_altpriority_encoder18_w_lg_zero239w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero237w238w(i);
	END GENERATE loop36;
	altpriority_encoder18 :  convert_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --convert_altpriority_encoder_r08

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END convert_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF convert_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero192w193w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero194w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero194w195w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  convert_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  convert_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero192w & wire_altpriority_encoder10_w_lg_w_lg_zero194w195w);
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero192w193w(i) <= wire_altpriority_encoder10_w_lg_zero192w(0) AND wire_altpriority_encoder10_q(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_zero194w(i) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(i);
	END GENERATE loop38;
	wire_altpriority_encoder10_w_lg_zero192w(0) <= NOT wire_altpriority_encoder10_zero;
	loop39 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero194w195w(i) <= wire_altpriority_encoder10_w_lg_zero194w(i) OR wire_altpriority_encoder10_w_lg_w_lg_zero192w193w(i);
	END GENERATE loop39;
	altpriority_encoder10 :  convert_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  convert_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --convert_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 1 reg 247 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  convert_altfp_convert_l1n IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END convert_altfp_convert_l1n;

 ARCHITECTURE RTL OF convert_altfp_convert_l1n IS

	 SIGNAL  wire_altbarrel_shift5_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 add_1_adder1_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q58w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_1_adder1_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_reg_w_lg_w_lg_q67w68w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q66w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissa_pre_round_reg_w_q_range59w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub6_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_w_lg_alb21w22w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb20w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cmpr4_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w52w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mantissa_overflow71w72w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector17w18w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow70w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector16w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range34w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range37w41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range40w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range43w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range46w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_adder1_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder2_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  mantissa_overflow :	STD_LOGIC;
	 SIGNAL  mantissa_post_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  sticky_bit_bus :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_or_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  convert_altbarrel_shift_tvf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  convert_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w(0) <= wire_w_lg_w_lg_guard_bit_w52w53w(0) AND sticky_bit_w;
	wire_w_lg_w_lg_guard_bit_w52w53w(0) <= wire_w_lg_guard_bit_w52w(0) AND round_bit_w;
	loop40 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_mantissa_overflow71w72w(i) <= wire_w_lg_mantissa_overflow71w(0) AND exponent_bus_pre_reg(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector17w18w(i) <= wire_w_lg_max_neg_value_selector17w(0) AND exponent_zero_w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_mantissa_overflow70w(i) <= mantissa_overflow AND wire_add_sub8_result(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_max_neg_value_selector16w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop45;
	wire_w_lg_guard_bit_w52w(0) <= NOT guard_bit_w;
	wire_w_lg_mantissa_overflow71w(0) <= NOT mantissa_overflow;
	wire_w_lg_max_neg_value_selector17w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	wire_w_lg_w_sticky_bit_or_w_range34w38w(0) <= wire_w_sticky_bit_or_w_range34w(0) OR wire_w_sticky_bit_bus_range36w(0);
	wire_w_lg_w_sticky_bit_or_w_range37w41w(0) <= wire_w_sticky_bit_or_w_range37w(0) OR wire_w_sticky_bit_bus_range39w(0);
	wire_w_lg_w_sticky_bit_or_w_range40w44w(0) <= wire_w_sticky_bit_or_w_range40w(0) OR wire_w_sticky_bit_bus_range42w(0);
	wire_w_lg_w_sticky_bit_or_w_range43w47w(0) <= wire_w_sticky_bit_or_w_range43w(0) OR wire_w_sticky_bit_bus_range45w(0);
	wire_w_lg_w_sticky_bit_or_w_range46w50w(0) <= wire_w_sticky_bit_or_w_range46w(0) OR wire_w_sticky_bit_bus_range48w(0);
	aclr <= '0';
	add_1_adder1_w <= add_1_adder1_reg;
	add_1_adder2_w <= (wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w OR wire_add_1_adder1_cout_reg_w_lg_q58w);
	add_1_adder_w <= ( add_1_adder2_w & add_1_adder1_w);
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w(0) OR (guard_bit_w AND round_bit_w));
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10011101";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector17w18w OR wire_w_lg_max_neg_value_selector16w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_cmpr4_w_lg_w_lg_alb21w22w OR wire_cmpr4_w_lg_alb20w);
	exponent_output_w <= wire_add_sub3_result;
	exponent_rounded <= (wire_w_lg_w_lg_mantissa_overflow71w72w OR wire_w_lg_mantissa_overflow70w);
	exponent_zero_w <= (OTHERS => '0');
	guard_bit_w <= shifted_mag_int_a(7);
	int_a <= dataa(30 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(22 DOWNTO 0);
	mantissa_overflow <= ((add_1_reg AND add_1_adder1_cout_reg) AND add_1_adder2_cout_reg);
	mantissa_post_round <= add_1_adder_w;
	mantissa_pre_round <= shifted_mag_int_a(30 DOWNTO 7);
	mantissa_rounded <= (wire_add_1_reg_w_lg_w_lg_q67w68w OR wire_add_1_reg_w_lg_q66w);
	max_neg_value_selector <= (wire_cmpr4_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10011110";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	round_bit_w <= shifted_mag_int_a(6);
	shifted_mag_int_a <= wire_altbarrel_shift5_result(30 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(31);
	sticky_bit_bus <= shifted_mag_int_a(5 DOWNTO 0);
	sticky_bit_or_w <= ( wire_w_lg_w_sticky_bit_or_w_range46w50w & wire_w_lg_w_sticky_bit_or_w_range43w47w & wire_w_lg_w_sticky_bit_or_w_range40w44w & wire_w_lg_w_sticky_bit_or_w_range37w41w & wire_w_lg_w_sticky_bit_or_w_range34w38w & sticky_bit_bus(0));
	sticky_bit_w <= sticky_bit_or_w(5);
	zero_padding_w <= (OTHERS => '0');
	wire_w_sticky_bit_bus_range36w(0) <= sticky_bit_bus(1);
	wire_w_sticky_bit_bus_range39w(0) <= sticky_bit_bus(2);
	wire_w_sticky_bit_bus_range42w(0) <= sticky_bit_bus(3);
	wire_w_sticky_bit_bus_range45w(0) <= sticky_bit_bus(4);
	wire_w_sticky_bit_bus_range48w(0) <= sticky_bit_bus(5);
	wire_w_sticky_bit_or_w_range34w(0) <= sticky_bit_or_w(0);
	wire_w_sticky_bit_or_w_range37w(0) <= sticky_bit_or_w(1);
	wire_w_sticky_bit_or_w_range40w(0) <= sticky_bit_or_w(2);
	wire_w_sticky_bit_or_w_range43w(0) <= sticky_bit_or_w(3);
	wire_w_sticky_bit_or_w_range46w(0) <= sticky_bit_or_w(4);
	wire_altbarrel_shift5_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift5 :  convert_altbarrel_shift_tvf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift5_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift5_result
	  );
	altpriority_encoder2 :  convert_altpriority_encoder_qb6
	  PORT MAP ( 
		data => prio_mag_int_a,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_cout_reg <= wire_add_sub6_cout;
			END IF;
		END IF;
	END PROCESS;
	loop46 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w(i) <= wire_add_1_adder1_cout_reg_w_lg_q60w(0) AND wire_mantissa_pre_round_reg_w_q_range59w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_q58w(i) <= add_1_adder1_cout_reg AND add_1_adder2_reg(i);
	END GENERATE loop47;
	wire_add_1_adder1_cout_reg_w_lg_q60w(0) <= NOT add_1_adder1_cout_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_reg <= wire_add_sub6_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_cout_reg <= wire_add_sub7_cout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_reg <= wire_add_sub7_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_reg <= add_1_w;
			END IF;
		END IF;
	END PROCESS;
	loop48 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_w_lg_q67w68w(i) <= wire_add_1_reg_w_lg_q67w(0) AND mantissa_pre_round_reg(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_q66w(i) <= add_1_reg AND mantissa_post_round(i);
	END GENERATE loop49;
	wire_add_1_reg_w_lg_q67w(0) <= NOT add_1_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	wire_mantissa_pre_round_reg_w_q_range59w <= mantissa_pre_round_reg(23 DOWNTO 12);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "0000000000000000000000000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 31,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_add_sub3_result
	  );
	wire_add_sub6_datab <= "000000000001";
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub6_cout,
		dataa => mantissa_pre_round(11 DOWNTO 0),
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	wire_add_sub7_datab <= "000000000001";
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub7_cout,
		dataa => mantissa_pre_round(23 DOWNTO 12),
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	wire_add_sub8_datab <= "00000001";
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_bus_pre_reg,
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	loop50 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_w_lg_alb21w22w(i) <= wire_cmpr4_w_lg_alb21w(0) AND exponent_output_w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_alb20w(i) <= wire_cmpr4_alb AND exceptions_value(i);
	END GENERATE loop51;
	wire_cmpr4_w_lg_alb21w(0) <= NOT wire_cmpr4_alb;
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr4_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --convert_altfp_convert_l1n
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY convert IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END convert;


ARCHITECTURE RTL OF convert IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT convert_altfp_convert_l1n
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	convert_altfp_convert_l1n_component : convert_altfp_convert_l1n
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "INT2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL convert.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: lpm
