-- megafunction wizard: %ALTFP_INV_SQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_INV_SQRT 

-- ============================================================
-- File Name: inv_sqrt.vhd
-- Megafunction Name(s):
-- 			ALTFP_INV_SQRT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_inv_sqrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=26 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altfp_inv_sqrt_and_or CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" LUT_INPUT_COUNT=4 OPERATION="OR" PIPELINE=3 WIDTH=23 aclr clken clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = reg 9 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_and_or_1de IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (22 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END inv_sqrt_altfp_inv_sqrt_and_or_1de;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_and_or_1de IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range378w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range406w410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range412w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range414w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range417w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range423w426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range425w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range428w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range381w385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range434w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range436w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range384w388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range390w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range392w396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range395w399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range401w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range403w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range450w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range453w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range456w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range462w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r3_w_range470w474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r3_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  operation_r3_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_connection_r2_w_range472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or5_w_operation_r3_w_range470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range378w382w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range378w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range380w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range406w410w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range406w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range408w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range412w415w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range412w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range413w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range414w418w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range414w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range416w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range417w421w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range417w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range419w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range423w426w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range423w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range424w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range425w429w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range425w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range427w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range428w432w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range428w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range430w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range381w385w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range381w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range383w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range434w437w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range434w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range435w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range436w440w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range436w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range438w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range384w388w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range384w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range386w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range390w393w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range390w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range391w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range392w396w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range392w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range394w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range395w399w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range395w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range397w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range401w404w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range401w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range402w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range403w407w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range403w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range405w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range450w454w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range450w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range452w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range453w457w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range453w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range455w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range456w460w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range456w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range458w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range462w465w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range462w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range463w(0);
	wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r3_w_range470w474w(0) <= wire_altfp_inv_sqrt_and_or5_w_operation_r3_w_range470w(0) OR wire_altfp_inv_sqrt_and_or5_w_connection_r2_w_range472w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	connection_r3_w <= connection_dffe2;
	operation_r1_w <= ( wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range436w440w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range434w437w & connection_r0_w(20) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range428w432w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range425w429w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range423w426w & connection_r0_w(16) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range417w421w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range414w418w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range412w415w & connection_r0_w(12) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range406w410w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range403w407w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range401w404w & connection_r0_w(8) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range395w399w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range392w396w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range390w393w & connection_r0_w(4) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range384w388w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range381w385w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r1_w_range378w382w & connection_r0_w(0));
	operation_r2_w <= ( wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range462w465w & connection_r1_w(4) & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range456w460w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range453w457w & wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r2_w_range450w454w & connection_r1_w(0));
	operation_r3_w <= ( wire_altfp_inv_sqrt_and_or5_w_lg_w_operation_r3_w_range470w474w & connection_r2_w(0));
	result <= connection_r3_w(0);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range405w(0) <= connection_r0_w(10);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range408w(0) <= connection_r0_w(11);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range413w(0) <= connection_r0_w(13);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range416w(0) <= connection_r0_w(14);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range419w(0) <= connection_r0_w(15);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range424w(0) <= connection_r0_w(17);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range427w(0) <= connection_r0_w(18);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range430w(0) <= connection_r0_w(19);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range380w(0) <= connection_r0_w(1);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range435w(0) <= connection_r0_w(21);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range438w(0) <= connection_r0_w(22);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range383w(0) <= connection_r0_w(2);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range386w(0) <= connection_r0_w(3);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range391w(0) <= connection_r0_w(5);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range394w(0) <= connection_r0_w(6);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range397w(0) <= connection_r0_w(7);
	wire_altfp_inv_sqrt_and_or5_w_connection_r0_w_range402w(0) <= connection_r0_w(9);
	wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range452w(0) <= connection_r1_w(1);
	wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range455w(0) <= connection_r1_w(2);
	wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range458w(0) <= connection_r1_w(3);
	wire_altfp_inv_sqrt_and_or5_w_connection_r1_w_range463w(0) <= connection_r1_w(5);
	wire_altfp_inv_sqrt_and_or5_w_connection_r2_w_range472w(0) <= connection_r2_w(1);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range378w(0) <= operation_r1_w(0);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range406w(0) <= operation_r1_w(10);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range412w(0) <= operation_r1_w(12);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range414w(0) <= operation_r1_w(13);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range417w(0) <= operation_r1_w(14);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range423w(0) <= operation_r1_w(16);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range425w(0) <= operation_r1_w(17);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range428w(0) <= operation_r1_w(18);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range381w(0) <= operation_r1_w(1);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range434w(0) <= operation_r1_w(20);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range436w(0) <= operation_r1_w(21);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range384w(0) <= operation_r1_w(2);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range390w(0) <= operation_r1_w(4);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range392w(0) <= operation_r1_w(5);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range395w(0) <= operation_r1_w(6);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range401w(0) <= operation_r1_w(8);
	wire_altfp_inv_sqrt_and_or5_w_operation_r1_w_range403w(0) <= operation_r1_w(9);
	wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range450w(0) <= operation_r2_w(0);
	wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range453w(0) <= operation_r2_w(1);
	wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range456w(0) <= operation_r2_w(2);
	wire_altfp_inv_sqrt_and_or5_w_operation_r2_w_range462w(0) <= operation_r2_w(4);
	wire_altfp_inv_sqrt_and_or5_w_operation_r3_w_range470w(0) <= operation_r3_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(22) & operation_r1_w(19) & operation_r1_w(15) & operation_r1_w(11) & operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1 <= ( operation_r2_w(5) & operation_r2_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2(0) <= ( operation_r3_w(1));
			END IF;
		END IF;
	END PROCESS;

 END RTL; --inv_sqrt_altfp_inv_sqrt_and_or_1de


--altfp_inv_sqrt_and_or CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" LUT_INPUT_COUNT=4 OPERATION="AND" PIPELINE=3 WIDTH=23 aclr clken clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = reg 9 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_and_or_jfe IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (22 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END inv_sqrt_altfp_inv_sqrt_and_or_jfe;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_and_or_jfe IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range479w483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range507w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range513w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range515w519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range518w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range524w527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range526w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range529w533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range482w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range535w538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range537w541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range485w489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range491w494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range493w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range496w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range502w505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range504w508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range551w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range554w558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range557w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range563w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r3_w_range571w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r3_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  operation_r3_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_connection_r2_w_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_w_operation_r3_w_range571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range479w483w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range479w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range481w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range507w511w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range507w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range509w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range513w516w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range513w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range514w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range515w519w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range515w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range517w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range518w522w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range518w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range520w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range524w527w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range524w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range525w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range526w530w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range526w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range528w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range529w533w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range529w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range531w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range482w486w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range482w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range484w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range535w538w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range535w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range536w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range537w541w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range537w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range539w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range485w489w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range485w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range487w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range491w494w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range491w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range492w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range493w497w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range493w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range495w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range496w500w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range496w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range498w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range502w505w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range502w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range503w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range504w508w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range504w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range506w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range551w555w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range551w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range553w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range554w558w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range554w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range556w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range557w561w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range557w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range559w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range563w566w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range563w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range564w(0);
	wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r3_w_range571w575w(0) <= wire_altfp_inv_sqrt_and_or6_w_operation_r3_w_range571w(0) AND wire_altfp_inv_sqrt_and_or6_w_connection_r2_w_range573w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	connection_r3_w <= connection_dffe2;
	operation_r1_w <= ( wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range537w541w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range535w538w & connection_r0_w(20) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range529w533w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range526w530w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range524w527w & connection_r0_w(16) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range518w522w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range515w519w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range513w516w & connection_r0_w(12) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range507w511w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range504w508w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range502w505w & connection_r0_w(8) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range496w500w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range493w497w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range491w494w & connection_r0_w(4) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range485w489w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range482w486w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r1_w_range479w483w & connection_r0_w(0));
	operation_r2_w <= ( wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range563w566w & connection_r1_w(4) & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range557w561w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range554w558w & wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r2_w_range551w555w & connection_r1_w(0));
	operation_r3_w <= ( wire_altfp_inv_sqrt_and_or6_w_lg_w_operation_r3_w_range571w575w & connection_r2_w(0));
	result <= connection_r3_w(0);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range506w(0) <= connection_r0_w(10);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range509w(0) <= connection_r0_w(11);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range514w(0) <= connection_r0_w(13);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range517w(0) <= connection_r0_w(14);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range520w(0) <= connection_r0_w(15);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range525w(0) <= connection_r0_w(17);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range528w(0) <= connection_r0_w(18);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range531w(0) <= connection_r0_w(19);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range481w(0) <= connection_r0_w(1);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range536w(0) <= connection_r0_w(21);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range539w(0) <= connection_r0_w(22);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range484w(0) <= connection_r0_w(2);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range487w(0) <= connection_r0_w(3);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range492w(0) <= connection_r0_w(5);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range495w(0) <= connection_r0_w(6);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range498w(0) <= connection_r0_w(7);
	wire_altfp_inv_sqrt_and_or6_w_connection_r0_w_range503w(0) <= connection_r0_w(9);
	wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range553w(0) <= connection_r1_w(1);
	wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range556w(0) <= connection_r1_w(2);
	wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range559w(0) <= connection_r1_w(3);
	wire_altfp_inv_sqrt_and_or6_w_connection_r1_w_range564w(0) <= connection_r1_w(5);
	wire_altfp_inv_sqrt_and_or6_w_connection_r2_w_range573w(0) <= connection_r2_w(1);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range479w(0) <= operation_r1_w(0);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range507w(0) <= operation_r1_w(10);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range513w(0) <= operation_r1_w(12);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range515w(0) <= operation_r1_w(13);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range518w(0) <= operation_r1_w(14);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range524w(0) <= operation_r1_w(16);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range526w(0) <= operation_r1_w(17);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range529w(0) <= operation_r1_w(18);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range482w(0) <= operation_r1_w(1);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range535w(0) <= operation_r1_w(20);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range537w(0) <= operation_r1_w(21);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range485w(0) <= operation_r1_w(2);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range491w(0) <= operation_r1_w(4);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range493w(0) <= operation_r1_w(5);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range496w(0) <= operation_r1_w(6);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range502w(0) <= operation_r1_w(8);
	wire_altfp_inv_sqrt_and_or6_w_operation_r1_w_range504w(0) <= operation_r1_w(9);
	wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range551w(0) <= operation_r2_w(0);
	wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range554w(0) <= operation_r2_w(1);
	wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range557w(0) <= operation_r2_w(2);
	wire_altfp_inv_sqrt_and_or6_w_operation_r2_w_range563w(0) <= operation_r2_w(4);
	wire_altfp_inv_sqrt_and_or6_w_operation_r3_w_range571w(0) <= operation_r3_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(22) & operation_r1_w(19) & operation_r1_w(15) & operation_r1_w(11) & operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1 <= ( operation_r2_w(5) & operation_r2_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2(0) <= ( operation_r3_w(1));
			END IF;
		END IF;
	END PROCESS;

 END RTL; --inv_sqrt_altfp_inv_sqrt_and_or_jfe


--altfp_inv_sqrt_and_or CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" LUT_INPUT_COUNT=4 OPERATION="OR" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_and_or_kbe IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END inv_sqrt_altfp_inv_sqrt_and_or_kbe;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_and_or_kbe IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range580w584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range583w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range586w590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range592w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range594w598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range597w601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r2_w_range607w611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_connection_r1_w_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_w_operation_r2_w_range607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range580w584w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range580w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range582w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range583w587w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range583w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range585w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range586w590w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range586w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range588w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range592w595w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range592w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range593w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range594w598w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range594w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range596w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range597w601w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range597w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range599w(0);
	wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r2_w_range607w611w(0) <= wire_altfp_inv_sqrt_and_or7_w_operation_r2_w_range607w(0) OR wire_altfp_inv_sqrt_and_or7_w_connection_r1_w_range609w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range597w601w & wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range594w598w & wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range592w595w & connection_r0_w(4) & wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range586w590w & wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range583w587w & wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r1_w_range580w584w & connection_r0_w(0));
	operation_r2_w <= ( wire_altfp_inv_sqrt_and_or7_w_lg_w_operation_r2_w_range607w611w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range582w(0) <= connection_r0_w(1);
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range585w(0) <= connection_r0_w(2);
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range588w(0) <= connection_r0_w(3);
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range593w(0) <= connection_r0_w(5);
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range596w(0) <= connection_r0_w(6);
	wire_altfp_inv_sqrt_and_or7_w_connection_r0_w_range599w(0) <= connection_r0_w(7);
	wire_altfp_inv_sqrt_and_or7_w_connection_r1_w_range609w(0) <= connection_r1_w(1);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range580w(0) <= operation_r1_w(0);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range583w(0) <= operation_r1_w(1);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range586w(0) <= operation_r1_w(2);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range592w(0) <= operation_r1_w(4);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range594w(0) <= operation_r1_w(5);
	wire_altfp_inv_sqrt_and_or7_w_operation_r1_w_range597w(0) <= operation_r1_w(6);
	wire_altfp_inv_sqrt_and_or7_w_operation_r2_w_range607w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --inv_sqrt_altfp_inv_sqrt_and_or_kbe


--altfp_inv_sqrt_and_or CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" LUT_INPUT_COUNT=4 OPERATION="AND" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_and_or_6ee IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END inv_sqrt_altfp_inv_sqrt_and_or_6ee;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_and_or_6ee IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range616w620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range619w623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range622w626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range628w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range630w634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range633w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r2_w_range643w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_connection_r1_w_range645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_w_operation_r2_w_range643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range616w620w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range616w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range618w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range619w623w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range619w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range621w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range622w626w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range622w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range624w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range628w631w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range628w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range629w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range630w634w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range630w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range632w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range633w637w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range633w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range635w(0);
	wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r2_w_range643w647w(0) <= wire_altfp_inv_sqrt_and_or8_w_operation_r2_w_range643w(0) AND wire_altfp_inv_sqrt_and_or8_w_connection_r1_w_range645w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range633w637w & wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range630w634w & wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range628w631w & connection_r0_w(4) & wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range622w626w & wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range619w623w & wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r1_w_range616w620w & connection_r0_w(0));
	operation_r2_w <= ( wire_altfp_inv_sqrt_and_or8_w_lg_w_operation_r2_w_range643w647w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range618w(0) <= connection_r0_w(1);
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range621w(0) <= connection_r0_w(2);
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range624w(0) <= connection_r0_w(3);
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range629w(0) <= connection_r0_w(5);
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range632w(0) <= connection_r0_w(6);
	wire_altfp_inv_sqrt_and_or8_w_connection_r0_w_range635w(0) <= connection_r0_w(7);
	wire_altfp_inv_sqrt_and_or8_w_connection_r1_w_range645w(0) <= connection_r1_w(1);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range616w(0) <= operation_r1_w(0);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range619w(0) <= operation_r1_w(1);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range622w(0) <= operation_r1_w(2);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range628w(0) <= operation_r1_w(4);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range630w(0) <= operation_r1_w(5);
	wire_altfp_inv_sqrt_and_or8_w_operation_r1_w_range633w(0) <= operation_r1_w(6);
	wire_altfp_inv_sqrt_and_or8_w_operation_r2_w_range643w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --inv_sqrt_altfp_inv_sqrt_and_or_6ee


--altfp_inv_sqrt_and_or CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" LUT_INPUT_COUNT=4 OPERATION="OR" PIPELINE=0 WIDTH=2 aclr clken clock data result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_and_or_bbe IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END inv_sqrt_altfp_inv_sqrt_and_or_bbe;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_and_or_bbe IS

	 SIGNAL  wire_stickybit_or0_w_lg_w_operation_r1_w_range652w656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stickybit_or0_w_connection_r0_w_range654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stickybit_or0_w_operation_r1_w_range652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_stickybit_or0_w_lg_w_operation_r1_w_range652w656w(0) <= wire_stickybit_or0_w_operation_r1_w_range652w(0) OR wire_stickybit_or0_w_connection_r0_w_range654w(0);
	connection_r0_w <= data;
	connection_r1_w(0) <= ( operation_r1_w(1));
	operation_r1_w <= ( wire_stickybit_or0_w_lg_w_operation_r1_w_range652w656w & connection_r0_w(0));
	result <= connection_r1_w(0);
	wire_stickybit_or0_w_connection_r0_w_range654w(0) <= connection_r0_w(1);
	wire_stickybit_or0_w_operation_r1_w_range652w(0) <= operation_r1_w(0);

 END RTL; --inv_sqrt_altfp_inv_sqrt_and_or_bbe


--altfp_inv_sqrt_csa CARRY_SELECT="YES" CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" DIRECTION="SUB" PIPELINE=1 REGISTER_INPUT="NO" REPRESENTATION="UNSIGNED" WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_csa_k4j IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END inv_sqrt_altfp_inv_sqrt_csa_k4j;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_csa_k4j IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout666w667w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout665w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout666w667w668w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  dataa_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  datab_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	dataa_w <= dataa;
	datab_w <= datab;
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout666w667w668w & wire_csa_lower_result);
	loop0 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout666w667w(i) <= wire_csa_lower_w_lg_cout666w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_cout665w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop1;
	wire_csa_lower_w_lg_cout666w(0) <= NOT wire_csa_lower_cout;
	loop2 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout666w667w668w(i) <= wire_csa_lower_w_lg_w_lg_cout666w667w(i) OR wire_csa_lower_w_lg_cout665w(i);
	END GENERATE loop2;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa_w(12 DOWNTO 0),
		datab => datab_w(12 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa_w(25 DOWNTO 13),
		datab => datab_w(25 DOWNTO 13),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa_w(25 DOWNTO 13),
		datab => datab_w(25 DOWNTO 13),
		result => wire_csa_upper1_result
	  );

 END RTL; --inv_sqrt_altfp_inv_sqrt_csa_k4j


--altfp_inv_sqrt_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" DIRECTION="ADD" PIPELINE=1 REGISTER_INPUT="NO" REPRESENTATION="UNSIGNED" WIDTH=13 aclr clken clock dataa datab result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_csa_rvi IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (12 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (12 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (12 DOWNTO 0)
	 ); 
 END inv_sqrt_altfp_inv_sqrt_csa_rvi;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_csa_rvi IS

	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  dataa_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  datab_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	dataa_w <= dataa;
	datab_w <= datab;
	result <= result_w;
	result_w <= wire_add_sub9_result;
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa_w,
		datab => datab_w,
		result => wire_add_sub9_result
	  );

 END RTL; --inv_sqrt_altfp_inv_sqrt_csa_rvi


--altfp_inv_sqrt_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" DIRECTION="SUB" PIPELINE=1 REGISTER_INPUT="NO" REPRESENTATION="UNSIGNED" WIDTH=13 aclr clken clock dataa datab result
--VERSION_BEGIN 13.0 cbx_altfp_inv_sqrt 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_mult 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_padd 2013:06:12:18:03:43:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_csa_s0j IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (12 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (12 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (12 DOWNTO 0)
	 ); 
 END inv_sqrt_altfp_inv_sqrt_csa_s0j;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_csa_s0j IS

	 SIGNAL  wire_add_sub10_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  dataa_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  datab_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	dataa_w <= dataa;
	datab_w <= datab;
	result <= result_w;
	result_w <= wire_add_sub10_result;
	add_sub10 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa_w,
		datab => datab_w,
		result => wire_add_sub10_result
	  );

 END RTL; --inv_sqrt_altfp_inv_sqrt_csa_s0j

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 16 lpm_mult 6 lpm_mux 1 reg 1094 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  inv_sqrt_altfp_inv_sqrt_s7d IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END inv_sqrt_altfp_inv_sqrt_s7d;

 ARCHITECTURE RTL OF inv_sqrt_altfp_inv_sqrt_s7d IS

	 SIGNAL  wire_altfp_inv_sqrt_and_or5_result	:	STD_LOGIC;
	 SIGNAL  wire_altfp_inv_sqrt_and_or6_result	:	STD_LOGIC;
	 SIGNAL  wire_altfp_inv_sqrt_and_or7_result	:	STD_LOGIC;
	 SIGNAL  wire_altfp_inv_sqrt_and_or8_result	:	STD_LOGIC;
	 SIGNAL  wire_stickybit_or0_result	:	STD_LOGIC;
	 SIGNAL  wire_stickybit_or1_result	:	STD_LOGIC;
	 SIGNAL  wire_diff_adder_0_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_diff_adder_1_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_slope_r1c1_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_slope_r1c2_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_slope_r1c3_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_slope_r2c1_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_slope_r2c2_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_slope_r3c1_add_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL	 and_dffe_0	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_dffe_1	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_dffe_2	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_dffe_3	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_dffe_4	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_dffe_5	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 division_by_zero_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_10	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_11	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_12	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_13	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_14	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_15	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_16	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_17	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_18	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_19	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_20	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_dffe1_20_w_lg_w_q_range325w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_dffe1_20_w_q_range325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exp_dffe1_3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_6	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_7	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_8	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe1_9	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe2_0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe2_1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe2_2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinite_input_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 intercept_dffe	:	STD_LOGIC_VECTOR(9 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_0	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_1	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_10	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_11	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_12	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_13	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_14	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_15	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_16	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_17	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_dffe_17_w_lg_w_lg_w_q_range272w276w277w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_dffe_17_w_lg_w_q_range272w274w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_dffe_17_w_lg_w_q_range272w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_dffe_17_w_q_range275w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_dffe_17_w_q_range273w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_man_dffe_17_w_q_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_dffe_2	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_3	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_4	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_5	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_6	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_7	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_8	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_dffe_9	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_input_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_output_dffe	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_dffe	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_0	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_1	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_10	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_11	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_12	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_13	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_2	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_3	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_4	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_5	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_6	:	STD_LOGIC_VECTOR(12 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_7	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_8	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_dffe_9	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_input_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_bias_adjustment_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_bias_adjustment_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_bias_adjustment_w_result_range342w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_inner_mult0_result	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_inner_mult1_result	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_outer_mult0_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_outer_mult1_result	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_sqr_mult0_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sqr_mult1_result	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_mux2_data_2d	:	STD_LOGIC_2D(47 DOWNTO 0, 15 DOWNTO 0);
	 SIGNAL  wire_mux2_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_mux2_w_result_range242w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_man_zero_w331w334w335w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_man_zero_w331w332w333w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_zero_w329w330w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_zero_w326w327w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_data_man_mux_w13w14w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinite_out_w365w366w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_zero_w331w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_zero_w331w332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_nan_input_w288w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_nan_out_w373w374w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_zero_out_w369w370w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_data_man_mux_w15w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinite_out_w367w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_zero_w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_zero_w326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_out_w375w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_out_w371w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range232w233w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range226w227w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range219w220w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range212w213w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range205w206w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_slope_w_range198w199w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_data_man_mux_w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_or_msb_w280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinite_out_w365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_or_msb_w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_zero_w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_input_w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_out_w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_out_w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  and_b0_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  and_b1_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  and_b2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  and_b3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  and_b4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  and_b5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  approx_c_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  approx_mx_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  approx_y_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  c_offset_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_3_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  const_bias_adj_eql_one_even_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  const_bias_adj_eql_one_odd_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  const_bias_adj_grt_one_even_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  const_bias_adj_grt_one_odd_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  const_bias_adj_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  data_exp_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  data_man_bus0_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  data_man_bus1_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  data_man_bus_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  data_man_mux_w :	STD_LOGIC;
	 SIGNAL  data_sign_w :	STD_LOGIC;
	 SIGNAL  division_by_zero_w :	STD_LOGIC;
	 SIGNAL  exp_and_msb_w :	STD_LOGIC;
	 SIGNAL  exp_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_exc_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_exc_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_one_w :	STD_LOGIC;
	 SIGNAL  exp_or_msb_w :	STD_LOGIC;
	 SIGNAL  exp_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_zero_w :	STD_LOGIC;
	 SIGNAL  gnd_w :	STD_LOGIC;
	 SIGNAL  infi_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  infinite_input_w :	STD_LOGIC;
	 SIGNAL  infinite_out_w :	STD_LOGIC;
	 SIGNAL  infinite_w :	STD_LOGIC;
	 SIGNAL  man_and_msb_w :	STD_LOGIC;
	 SIGNAL  man_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_exc_nan_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_exc_zeros_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_non_zero_w :	STD_LOGIC;
	 SIGNAL  man_one_w :	STD_LOGIC;
	 SIGNAL  man_or_msb_w :	STD_LOGIC;
	 SIGNAL  man_out_0_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_out_1_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_out_round_0_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_out_round_1_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_res_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_zero_w :	STD_LOGIC;
	 SIGNAL  modified_c_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  mux_1_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mux_2_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mux_3_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  nan_input_w :	STD_LOGIC;
	 SIGNAL  nan_out_w :	STD_LOGIC;
	 SIGNAL  nan_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  nan_w :	STD_LOGIC;
	 SIGNAL  norm_res_int_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  selector_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  shift_b0_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shift_b1_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shift_b2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shift_b3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shift_b4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shift_b5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sign_exc_bit_w :	STD_LOGIC;
	 SIGNAL  sign_res_w :	STD_LOGIC;
	 SIGNAL  slope_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  table_bus_full_w :	STD_LOGIC_VECTOR (767 DOWNTO 0);
	 SIGNAL  vcc_w :	STD_LOGIC;
	 SIGNAL  x_0_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  x_1_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  x_2_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  x_initial_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  zero_input_w :	STD_LOGIC;
	 SIGNAL  zero_one_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  zero_out_w :	STD_LOGIC;
	 SIGNAL  zero_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  zero_w :	STD_LOGIC;
	 SIGNAL  wire_w_and_b0_w_range200w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_and_b1_w_range207w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_and_b2_w_range214w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_and_b3_w_range221w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_and_b4_w_range228w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_and_b5_w_range234w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_slope_w_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_and_or_1de
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_and_or_jfe
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_and_or_kbe
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_and_or_6ee
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_and_or_bbe
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_csa_k4j
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_csa_rvi
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(12 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(12 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(12 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  inv_sqrt_altfp_inv_sqrt_csa_s0j
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(12 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(12 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(12 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop3 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_man_zero_w331w334w335w(i) <= wire_w_lg_w_lg_man_zero_w331w334w(0) AND const_bias_adj_grt_one_even_w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_man_zero_w331w332w333w(i) <= wire_w_lg_w_lg_man_zero_w331w332w(0) AND const_bias_adj_grt_one_odd_w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_man_zero_w329w330w(i) <= wire_w_lg_man_zero_w329w(0) AND const_bias_adj_eql_one_even_w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_man_zero_w326w327w(i) <= wire_w_lg_man_zero_w326w(0) AND const_bias_adj_eql_one_odd_w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_w_lg_data_man_mux_w13w14w(i) <= wire_w_lg_data_man_mux_w13w(0) AND data_man_bus1_w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_infinite_out_w365w366w(i) <= wire_w_lg_infinite_out_w365w(0) AND norm_res_int_w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_man_zero_w331w334w(0) <= wire_w_lg_man_zero_w331w(0) AND wire_exp_dffe1_20_w_lg_w_q_range325w328w(0);
	wire_w_lg_w_lg_man_zero_w331w332w(0) <= wire_w_lg_man_zero_w331w(0) AND wire_exp_dffe1_20_w_q_range325w(0);
	wire_w_lg_w_lg_nan_input_w288w289w(0) <= wire_w_lg_nan_input_w288w(0) AND infinite_input_w;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_nan_out_w373w374w(i) <= wire_w_lg_nan_out_w373w(0) AND mux_2_res_w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_zero_out_w369w370w(i) <= wire_w_lg_zero_out_w369w(0) AND mux_1_res_w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_data_man_mux_w15w(i) <= data_man_mux_w AND data_man_bus0_w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_infinite_out_w367w(i) <= infinite_out_w AND infi_res_w(i);
	END GENERATE loop12;
	wire_w_lg_man_zero_w329w(0) <= man_zero_w AND wire_exp_dffe1_20_w_lg_w_q_range325w328w(0);
	wire_w_lg_man_zero_w326w(0) <= man_zero_w AND wire_exp_dffe1_20_w_q_range325w(0);
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_nan_out_w375w(i) <= nan_out_w AND nan_res_w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_zero_out_w371w(i) <= zero_out_w AND zero_res_w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range232w233w(i) <= wire_w_slope_w_range232w(0) AND shift_b5_w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range226w227w(i) <= wire_w_slope_w_range226w(0) AND shift_b4_w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range219w220w(i) <= wire_w_slope_w_range219w(0) AND shift_b3_w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range212w213w(i) <= wire_w_slope_w_range212w(0) AND shift_b2_w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range205w206w(i) <= wire_w_slope_w_range205w(0) AND shift_b1_w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_slope_w_range198w199w(i) <= wire_w_slope_w_range198w(0) AND shift_b0_w(i);
	END GENERATE loop20;
	wire_w_lg_data_man_mux_w13w(0) <= NOT data_man_mux_w;
	wire_w_lg_exp_or_msb_w280w(0) <= NOT exp_or_msb_w;
	wire_w_lg_infinite_out_w365w(0) <= NOT infinite_out_w;
	wire_w_lg_man_or_msb_w279w(0) <= NOT man_or_msb_w;
	wire_w_lg_man_zero_w331w(0) <= NOT man_zero_w;
	wire_w_lg_nan_input_w288w(0) <= NOT nan_input_w;
	wire_w_lg_nan_out_w373w(0) <= NOT nan_out_w;
	wire_w_lg_zero_out_w369w(0) <= NOT zero_out_w;
	aclr <= '0';
	and_b0_w <= wire_w_lg_w_slope_w_range198w199w;
	and_b1_w <= wire_w_lg_w_slope_w_range205w206w;
	and_b2_w <= wire_w_lg_w_slope_w_range212w213w;
	and_b3_w <= wire_w_lg_w_slope_w_range219w220w;
	and_b4_w <= wire_w_lg_w_slope_w_range226w227w;
	and_b5_w <= wire_w_lg_w_slope_w_range232w233w;
	approx_c_w <= "1110001";
	approx_mx_w <= ( gnd_w & man_dffe_0(24 DOWNTO 19));
	approx_y_w <= ( wire_add_sub3_result & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w);
	c_offset_w <= ( gnd_w & gnd_w & gnd_w & intercept_dffe);
	clk_en <= '1';
	const_3_w <= "11000000000000000000000000";
	const_bias_adj_eql_one_even_w <= "101111100";
	const_bias_adj_eql_one_odd_w <= "101111101";
	const_bias_adj_grt_one_even_w <= "101111100";
	const_bias_adj_grt_one_odd_w <= "101111011";
	const_bias_adj_w <= (((wire_w_lg_w_lg_w_lg_man_zero_w331w334w335w OR wire_w_lg_w_lg_w_lg_man_zero_w331w332w333w) OR wire_w_lg_w_lg_man_zero_w329w330w) OR wire_w_lg_w_lg_man_zero_w326w327w);
	data_exp_bus_w <= data(30 DOWNTO 23);
	data_man_bus0_w <= ( gnd_w & vcc_w & data(22 DOWNTO 0));
	data_man_bus1_w <= ( vcc_w & data(22 DOWNTO 0) & gnd_w);
	data_man_bus_w <= (wire_w_lg_data_man_mux_w15w OR wire_w_lg_w_lg_data_man_mux_w13w14w);
	data_man_mux_w <= data(23);
	data_sign_w <= data(31);
	division_by_zero_w <= (zero_input_w AND (NOT sign_dffe(21)));
	exp_and_msb_w <= wire_altfp_inv_sqrt_and_or8_result;
	exp_bus_w <= exp_dffe1_17;
	exp_exc_ones_w <= (OTHERS => '1');
	exp_exc_zeros_w <= (OTHERS => '0');
	exp_one_w <= exp_and_msb_w;
	exp_or_msb_w <= wire_altfp_inv_sqrt_and_or7_result;
	exp_res_w <= exp_dffe2_2;
	exp_zero_w <= wire_w_lg_exp_or_msb_w280w(0);
	gnd_w <= '0';
	infi_res_w <= ( sign_exc_bit_w & exp_exc_ones_w & man_exc_zeros_w);
	infinite_input_w <= infinite_input_dffe;
	infinite_out_w <= infinite_dffe(2);
	infinite_w <= zero_input_w;
	man_and_msb_w <= wire_altfp_inv_sqrt_and_or6_result;
	man_bus_w <= (wire_man_dffe_17_w_lg_w_lg_w_q_range272w276w277w OR wire_man_dffe_17_w_lg_w_q_range272w274w);
	man_exc_nan_w <= ( vcc_w & man_exc_zeros_w(21 DOWNTO 0));
	man_exc_zeros_w <= (OTHERS => '0');
	man_non_zero_w <= man_or_msb_w;
	man_one_w <= man_and_msb_w;
	man_or_msb_w <= wire_altfp_inv_sqrt_and_or5_result;
	man_out_0_w <= man_out_round_0_w;
	man_out_1_w <= man_out_round_1_w;
	man_out_round_0_w <= ( man_dffe_7(24 DOWNTO 2) & wire_stickybit_or0_result);
	man_out_round_1_w <= ( man_dffe_17(24 DOWNTO 2) & wire_stickybit_or1_result);
	man_res_w <= x_2_w(22 DOWNTO 0);
	man_zero_w <= wire_w_lg_man_or_msb_w279w(0);
	modified_c_w <= wire_add_sub4_result(12 DOWNTO 0);
	mux_1_res_w <= (wire_w_lg_infinite_out_w367w OR wire_w_lg_w_lg_infinite_out_w365w366w);
	mux_2_res_w <= (wire_w_lg_zero_out_w371w OR wire_w_lg_w_lg_zero_out_w369w370w);
	mux_3_res_w <= (wire_w_lg_nan_out_w375w OR wire_w_lg_w_lg_nan_out_w373w374w);
	nan_input_w <= nan_input_dffe;
	nan_out_w <= nan_dffe(2);
	nan_res_w <= ( sign_exc_bit_w & exp_exc_ones_w & man_exc_nan_w);
	nan_w <= (nan_input_w OR sign_dffe(21));
	norm_res_int_w <= ( sign_res_w & exp_res_w & man_res_w);
	result <= result_output_dffe;
	selector_w <= ( wire_add_sub1_result & data_man_bus_w(22 DOWNTO 19));
	shift_b0_w <= ( gnd_w & gnd_w & man_dffe_0 & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w);
	shift_b1_w <= ( gnd_w & gnd_w & gnd_w & man_dffe_0 & gnd_w & gnd_w & gnd_w & gnd_w);
	shift_b2_w <= ( gnd_w & gnd_w & gnd_w & gnd_w & man_dffe_0 & gnd_w & gnd_w & gnd_w);
	shift_b3_w <= ( gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & man_dffe_0 & gnd_w & gnd_w);
	shift_b4_w <= ( gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & man_dffe_0 & gnd_w);
	shift_b5_w <= ( gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & gnd_w & man_dffe_0);
	sign_exc_bit_w <= sign_res_w;
	sign_res_w <= sign_dffe(24);
	slope_w <= wire_mux2_result(15 DOWNTO 10);
	table_bus_full_w <= ( "0010010000000011" & "0010010001000100" & "0010010010000100" & "0010010011000100" & "0010010100000100" & "0010100011010001" & "0010100100010010" & "0010100101010010" & "0010100110010010" & "0010110101100111" & "0010110110100111" & "0010110111100111" & "0011000111000010" & "0011001000000011" & "0011001001000011" & "0011011000100011" & "0011011001100100" & "0011011010100100" & "0011101010001001" & "0011101011001010" & "0011111010110011" & "0011111011110011" & "0100001011100001" & "0100001100100001" & "0100011100010010" & "0100101100000110" & "0100101101000110" & "0100111100111101" & "0101001100110110" & "0101011100110010" & "0101101100101111" & "0101111100101111" & "0110001100110001" & "0110011100110100" & "0110101100111001" & "0110111100111111" & "0111011100010000" & "0111111011100110" & "1000001011110011" & "1000101011001111" & "1001001010101111" & "1001111001100111" & "1010101000100100" & "1011010111101000" & "1100000110110001" & "1101000101011010" & "1110000100001010" & "1111100010000000");
	vcc_w <= '1';
	x_0_w <= x_initial_w;
	x_1_w <= ( gnd_w & wire_outer_mult0_result(36 DOWNTO 13));
	x_2_w <= ( gnd_w & wire_outer_mult1_result(48 DOWNTO 25));
	x_initial_w <= wire_slope_r3c1_add_result;
	zero_input_w <= zero_input_dffe;
	zero_one_w <= "01";
	zero_out_w <= zero_dffe(2);
	zero_res_w <= ( sign_exc_bit_w & exp_exc_zeros_w & man_exc_zeros_w);
	zero_w <= (wire_w_lg_w_lg_nan_input_w288w289w(0) AND (NOT sign_dffe(21)));
	wire_w_and_b0_w_range200w <= and_b0_w(30 DOWNTO 18);
	wire_w_and_b1_w_range207w <= and_b1_w(30 DOWNTO 18);
	wire_w_and_b2_w_range214w <= and_b2_w(30 DOWNTO 18);
	wire_w_and_b3_w_range221w <= and_b3_w(30 DOWNTO 18);
	wire_w_and_b4_w_range228w <= and_b4_w(30 DOWNTO 18);
	wire_w_and_b5_w_range234w <= and_b5_w(30 DOWNTO 18);
	wire_w_slope_w_range232w(0) <= slope_w(0);
	wire_w_slope_w_range226w(0) <= slope_w(1);
	wire_w_slope_w_range219w(0) <= slope_w(2);
	wire_w_slope_w_range212w(0) <= slope_w(3);
	wire_w_slope_w_range205w(0) <= slope_w(4);
	wire_w_slope_w_range198w(0) <= slope_w(5);
	altfp_inv_sqrt_and_or5 :  inv_sqrt_altfp_inv_sqrt_and_or_1de
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_bus_w,
		result => wire_altfp_inv_sqrt_and_or5_result
	  );
	altfp_inv_sqrt_and_or6 :  inv_sqrt_altfp_inv_sqrt_and_or_jfe
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_bus_w,
		result => wire_altfp_inv_sqrt_and_or6_result
	  );
	altfp_inv_sqrt_and_or7 :  inv_sqrt_altfp_inv_sqrt_and_or_kbe
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_bus_w,
		result => wire_altfp_inv_sqrt_and_or7_result
	  );
	altfp_inv_sqrt_and_or8 :  inv_sqrt_altfp_inv_sqrt_and_or_6ee
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_bus_w,
		result => wire_altfp_inv_sqrt_and_or8_result
	  );
	stickybit_or0 :  inv_sqrt_altfp_inv_sqrt_and_or_bbe
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_dffe_7(1 DOWNTO 0),
		result => wire_stickybit_or0_result
	  );
	stickybit_or1 :  inv_sqrt_altfp_inv_sqrt_and_or_bbe
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_dffe_17(1 DOWNTO 0),
		result => wire_stickybit_or1_result
	  );
	diff_adder_0 :  inv_sqrt_altfp_inv_sqrt_csa_k4j
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => const_3_w(25 DOWNTO 0),
		datab => wire_inner_mult0_result(47 DOWNTO 22),
		result => wire_diff_adder_0_result
	  );
	diff_adder_1 :  inv_sqrt_altfp_inv_sqrt_csa_k4j
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => const_3_w(25 DOWNTO 0),
		datab => wire_inner_mult1_result(47 DOWNTO 22),
		result => wire_diff_adder_1_result
	  );
	slope_r1c1_add :  inv_sqrt_altfp_inv_sqrt_csa_rvi
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => and_dffe_0,
		datab => and_dffe_1,
		result => wire_slope_r1c1_add_result
	  );
	slope_r1c2_add :  inv_sqrt_altfp_inv_sqrt_csa_rvi
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => and_dffe_2,
		datab => and_dffe_3,
		result => wire_slope_r1c2_add_result
	  );
	slope_r1c3_add :  inv_sqrt_altfp_inv_sqrt_csa_rvi
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => and_dffe_4,
		datab => and_dffe_5,
		result => wire_slope_r1c3_add_result
	  );
	slope_r2c1_add :  inv_sqrt_altfp_inv_sqrt_csa_rvi
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_slope_r1c1_add_result,
		datab => wire_slope_r1c2_add_result,
		result => wire_slope_r2c1_add_result
	  );
	slope_r2c2_add :  inv_sqrt_altfp_inv_sqrt_csa_s0j
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => modified_c_w,
		datab => wire_slope_r1c3_add_result,
		result => wire_slope_r2c2_add_result
	  );
	slope_r3c1_add :  inv_sqrt_altfp_inv_sqrt_csa_s0j
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_slope_r2c2_add_result,
		datab => wire_slope_r2c1_add_result,
		result => wire_slope_r3c1_add_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_0 <= wire_w_and_b0_w_range200w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_1 <= wire_w_and_b1_w_range207w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_2 <= wire_w_and_b2_w_range214w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_3 <= wire_w_and_b3_w_range221w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_4 <= wire_w_and_b4_w_range228w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_dffe_5 <= wire_w_and_b5_w_range234w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN division_by_zero_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN division_by_zero_dffe <= ( division_by_zero_dffe(1 DOWNTO 0) & division_by_zero_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_0 <= data_exp_bus_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_1 <= exp_dffe1_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_10 <= exp_dffe1_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_11 <= exp_dffe1_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_12 <= exp_dffe1_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_13 <= exp_dffe1_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_14 <= exp_dffe1_13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_15 <= exp_dffe1_14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_16 <= exp_dffe1_15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_17 <= exp_dffe1_16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_18 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_18 <= exp_dffe1_17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_19 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_19 <= exp_dffe1_18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_2 <= exp_dffe1_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_20 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_20 <= exp_dffe1_19;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_dffe1_20_w_lg_w_q_range325w328w(0) <= NOT wire_exp_dffe1_20_w_q_range325w(0);
	wire_exp_dffe1_20_w_q_range325w(0) <= exp_dffe1_20(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_3 <= exp_dffe1_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_4 <= exp_dffe1_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_5 <= exp_dffe1_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_6 <= exp_dffe1_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_7 <= exp_dffe1_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_8 <= exp_dffe1_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1_9 <= exp_dffe1_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe2_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe2_0 <= wire_bias_adjustment_w_result_range342w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe2_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe2_1 <= exp_dffe2_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe2_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe2_2 <= exp_dffe2_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_dffe <= ( infinite_dffe(1 DOWNTO 0) & infinite_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinite_input_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinite_input_dffe <= (exp_one_w AND man_zero_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN intercept_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN intercept_dffe <= wire_mux2_w_result_range242w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_0 <= data_man_bus_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_1 <= man_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_10 <= man_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_11 <= man_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_12 <= man_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_13 <= man_dffe_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_14 <= man_dffe_13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_15 <= man_dffe_14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_16 <= man_dffe_15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_17 <= man_dffe_16;
			END IF;
		END IF;
	END PROCESS;
	loop21 : FOR i IN 0 TO 22 GENERATE 
		wire_man_dffe_17_w_lg_w_lg_w_q_range272w276w277w(i) <= wire_man_dffe_17_w_lg_w_q_range272w276w(0) AND wire_man_dffe_17_w_q_range275w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 22 GENERATE 
		wire_man_dffe_17_w_lg_w_q_range272w274w(i) <= wire_man_dffe_17_w_q_range272w(0) AND wire_man_dffe_17_w_q_range273w(i);
	END GENERATE loop22;
	wire_man_dffe_17_w_lg_w_q_range272w276w(0) <= NOT wire_man_dffe_17_w_q_range272w(0);
	wire_man_dffe_17_w_q_range275w <= man_dffe_17(22 DOWNTO 0);
	wire_man_dffe_17_w_q_range273w <= man_dffe_17(23 DOWNTO 1);
	wire_man_dffe_17_w_q_range272w(0) <= man_dffe_17(24);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_2 <= man_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_3 <= man_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_4 <= man_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_5 <= man_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_6 <= man_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_7 <= man_dffe_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_8 <= man_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_dffe_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_dffe_9 <= man_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_dffe <= ( nan_dffe(1 DOWNTO 0) & nan_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_input_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_input_dffe <= (exp_one_w AND (man_non_zero_w OR man_one_w));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_output_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_output_dffe <= mux_3_res_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_dffe <= ( sign_dffe(23 DOWNTO 0) & data_sign_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_0 <= x_0_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_1 <= x_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_10 <= x_dffe_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_11 <= x_dffe_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_12 <= x_dffe_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_13 <= x_dffe_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_2 <= x_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_3 <= x_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_4 <= x_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_5 <= x_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_6 <= x_dffe_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_7 <= x_1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_8 <= x_dffe_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_dffe_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN x_dffe_9 <= x_dffe_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_dffe <= ( zero_dffe(1 DOWNTO 0) & zero_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_input_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_input_dffe <= (exp_zero_w AND ((man_one_w OR man_non_zero_w) OR man_zero_w));
			END IF;
		END IF;
	END PROCESS;
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 2
	  )
	  PORT MAP ( 
		dataa => data_man_bus_w(24 DOWNTO 23),
		datab => zero_one_w,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => approx_c_w,
		datab => approx_mx_w,
		result => wire_add_sub3_result
	  );
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => approx_y_w,
		datab => c_offset_w,
		result => wire_add_sub4_result
	  );
	wire_bias_adjustment_datab <= ( gnd_w & exp_dffe1_20);
	wire_bias_adjustment_w_result_range342w <= wire_bias_adjustment_result(8 DOWNTO 1);
	bias_adjustment :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => const_bias_adj_w,
		datab => wire_bias_adjustment_datab,
		result => wire_bias_adjustment_result
	  );
	inner_mult0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 24,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 49,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_out_0_w,
		datab => wire_sqr_mult0_result(24 DOWNTO 0),
		result => wire_inner_mult0_result
	  );
	inner_mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 24,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 49,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_out_1_w,
		datab => wire_sqr_mult1_result(48 DOWNTO 24),
		result => wire_inner_mult1_result
	  );
	outer_mult0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 26,
		LPM_WIDTHB => 13,
		LPM_WIDTHP => 39,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_diff_adder_0_result(25 DOWNTO 0),
		datab => x_dffe_6,
		result => wire_outer_mult0_result
	  );
	outer_mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 26,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 51,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_diff_adder_1_result(25 DOWNTO 0),
		datab => x_dffe_13,
		result => wire_outer_mult1_result
	  );
	sqr_mult0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 13,
		LPM_WIDTHB => 13,
		LPM_WIDTHP => 26,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => x_0_w,
		datab => x_0_w,
		result => wire_sqr_mult0_result
	  );
	sqr_mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 25,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 50,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=AUTO"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => x_1_w,
		datab => x_1_w,
		result => wire_sqr_mult1_result
	  );
	loop23 : FOR i IN 0 TO 47 GENERATE
		loop24 : FOR j IN 0 TO 15 GENERATE
			wire_mux2_data_2d(i, j) <= table_bus_full_w(i*16+j);
		END GENERATE loop24;
	END GENERATE loop23;
	wire_mux2_w_result_range242w <= wire_mux2_result(9 DOWNTO 0);
	mux2 :  lpm_mux
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_SIZE => 48,
		LPM_WIDTH => 16,
		LPM_WIDTHS => 6
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => wire_mux2_data_2d,
		result => wire_mux2_result,
		sel => selector_w
	  );

 END RTL; --inv_sqrt_altfp_inv_sqrt_s7d
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY inv_sqrt IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END inv_sqrt;


ARCHITECTURE RTL OF inv_sqrt IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT inv_sqrt_altfp_inv_sqrt_s7d
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	inv_sqrt_altfp_inv_sqrt_s7d_component : inv_sqrt_altfp_inv_sqrt_s7d
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_inv_sqrt"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "26"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL inv_sqrt.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: lpm
