-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: converter.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" OPERATION="FLOAT2INT" ROUNDING="TO_NEAREST" WIDTH_DATA=32 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=9 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=9 clock dataa result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_altfp_convert 2013:06:12:18:03:43:SJ cbx_altpriority_encoder 2013:06:12:18:03:43:SJ cbx_altsyncram 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_abs 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_decode 2013:06:12:18:03:43:SJ cbx_lpm_divide 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_stratixiii 2013:06:12:18:03:43:SJ cbx_stratixv 2013:06:12:18:03:43:SJ cbx_util_mgl 2013:06:12:18:03:43:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=31 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ  VERSION_END

--synthesis_resources = reg 66 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  converter_altbarrel_shift_svf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (30 DOWNTO 0)
	 ); 
 END converter_altbarrel_shift_svf;

 ARCHITECTURE RTL OF converter_altbarrel_shift_svf IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w299w300w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w295w296w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w320w321w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w316w317w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w342w343w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w338w339w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w364w365w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w360w361w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w383w384w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w379w380w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w291w292w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w312w313w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w334w335w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w356w357w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w375w376w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range286w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range286w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range307w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range307w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range329w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range329w338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range352w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range352w360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range371w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range371w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range283w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range305w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range326w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range350w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_dir_w_range369w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range286w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range307w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range329w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range352w356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_sel_w_range371w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range286w299w300w301w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range307w320w321w322w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range329w342w343w344w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range352w364w365w366w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range371w383w384w385w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w302w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w323w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w345w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w367w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w386w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (185 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (154 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w294w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w297w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w315w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w318w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w337w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w340w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w359w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w362w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w378w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w381w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_dir_w_range369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range346w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range368w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range281w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range304w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sbit_w_range324w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_sel_w_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_smux_w_range374w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift6_w_smux_w_range333w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w299w300w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range286w299w(0) AND wire_altbarrel_shift6_w297w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w295w296w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range286w295w(0) AND wire_altbarrel_shift6_w294w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w320w321w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range307w320w(0) AND wire_altbarrel_shift6_w318w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w316w317w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range307w316w(0) AND wire_altbarrel_shift6_w315w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w342w343w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range329w342w(0) AND wire_altbarrel_shift6_w340w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w338w339w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range329w338w(0) AND wire_altbarrel_shift6_w337w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w364w365w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range352w364w(0) AND wire_altbarrel_shift6_w362w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w360w361w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range352w360w(0) AND wire_altbarrel_shift6_w359w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w383w384w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range371w383w(0) AND wire_altbarrel_shift6_w381w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w379w380w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range371w379w(0) AND wire_altbarrel_shift6_w378w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w291w292w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range286w291w(0) AND wire_altbarrel_shift6_w_sbit_w_range281w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w312w313w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range307w312w(0) AND wire_altbarrel_shift6_w_sbit_w_range304w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w334w335w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range329w334w(0) AND wire_altbarrel_shift6_w_sbit_w_range324w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w356w357w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range352w356w(0) AND wire_altbarrel_shift6_w_sbit_w_range346w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w375w376w(i) <= wire_altbarrel_shift6_w_lg_w_sel_w_range371w375w(0) AND wire_altbarrel_shift6_w_sbit_w_range368w(i);
	END GENERATE loop14;
	wire_altbarrel_shift6_w_lg_w_sel_w_range286w299w(0) <= wire_altbarrel_shift6_w_sel_w_range286w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range283w298w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range286w295w(0) <= wire_altbarrel_shift6_w_sel_w_range286w(0) AND wire_altbarrel_shift6_w_dir_w_range283w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range307w320w(0) <= wire_altbarrel_shift6_w_sel_w_range307w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range305w319w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range307w316w(0) <= wire_altbarrel_shift6_w_sel_w_range307w(0) AND wire_altbarrel_shift6_w_dir_w_range305w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range329w342w(0) <= wire_altbarrel_shift6_w_sel_w_range329w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range326w341w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range329w338w(0) <= wire_altbarrel_shift6_w_sel_w_range329w(0) AND wire_altbarrel_shift6_w_dir_w_range326w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range352w364w(0) <= wire_altbarrel_shift6_w_sel_w_range352w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range350w363w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range352w360w(0) <= wire_altbarrel_shift6_w_sel_w_range352w(0) AND wire_altbarrel_shift6_w_dir_w_range350w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range371w383w(0) <= wire_altbarrel_shift6_w_sel_w_range371w(0) AND wire_altbarrel_shift6_w_lg_w_dir_w_range369w382w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range371w379w(0) <= wire_altbarrel_shift6_w_sel_w_range371w(0) AND wire_altbarrel_shift6_w_dir_w_range369w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range283w298w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range283w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range305w319w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range305w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range326w341w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range326w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range350w363w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range350w(0);
	wire_altbarrel_shift6_w_lg_w_dir_w_range369w382w(0) <= NOT wire_altbarrel_shift6_w_dir_w_range369w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range286w291w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range286w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range307w312w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range307w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range329w334w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range329w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range352w356w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range352w(0);
	wire_altbarrel_shift6_w_lg_w_sel_w_range371w375w(0) <= NOT wire_altbarrel_shift6_w_sel_w_range371w(0);
	loop15 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range286w299w300w301w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w299w300w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w295w296w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range307w320w321w322w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w320w321w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w316w317w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range329w342w343w344w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w342w343w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w338w339w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range352w364w365w366w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w364w365w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w360w361w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range371w383w384w385w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w383w384w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w379w380w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w302w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range286w299w300w301w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range286w291w292w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w323w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range307w320w321w322w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range307w312w313w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w345w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range329w342w343w344w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range329w334w335w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w367w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range352w364w365w366w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range352w356w357w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 30 GENERATE 
		wire_altbarrel_shift6_w386w(i) <= wire_altbarrel_shift6_w_lg_w_lg_w_lg_w_sel_w_range371w383w384w385w(i) OR wire_altbarrel_shift6_w_lg_w_lg_w_sel_w_range371w375w376w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(1) & dir_w(3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(185 DOWNTO 155);
	sbit_w <= ( sbit_piper2d & smux_w(123 DOWNTO 93) & sbit_piper1d & smux_w(61 DOWNTO 0) & data);
	sel_w <= ( sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift6_w386w & wire_altbarrel_shift6_w367w & wire_altbarrel_shift6_w345w & wire_altbarrel_shift6_w323w & wire_altbarrel_shift6_w302w);
	wire_altbarrel_shift6_w294w <= ( pad_w(0) & sbit_w(30 DOWNTO 1));
	wire_altbarrel_shift6_w297w <= ( sbit_w(29 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift6_w315w <= ( pad_w(1 DOWNTO 0) & sbit_w(61 DOWNTO 33));
	wire_altbarrel_shift6_w318w <= ( sbit_w(59 DOWNTO 31) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift6_w337w <= ( pad_w(3 DOWNTO 0) & sbit_w(92 DOWNTO 66));
	wire_altbarrel_shift6_w340w <= ( sbit_w(88 DOWNTO 62) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift6_w359w <= ( pad_w(7 DOWNTO 0) & sbit_w(123 DOWNTO 101));
	wire_altbarrel_shift6_w362w <= ( sbit_w(115 DOWNTO 93) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift6_w378w <= ( pad_w(15 DOWNTO 0) & sbit_w(154 DOWNTO 140));
	wire_altbarrel_shift6_w381w <= ( sbit_w(138 DOWNTO 124) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift6_w_dir_w_range283w(0) <= dir_w(0);
	wire_altbarrel_shift6_w_dir_w_range305w(0) <= dir_w(1);
	wire_altbarrel_shift6_w_dir_w_range326w(0) <= dir_w(2);
	wire_altbarrel_shift6_w_dir_w_range350w(0) <= dir_w(3);
	wire_altbarrel_shift6_w_dir_w_range369w(0) <= dir_w(4);
	wire_altbarrel_shift6_w_sbit_w_range346w <= sbit_w(123 DOWNTO 93);
	wire_altbarrel_shift6_w_sbit_w_range368w <= sbit_w(154 DOWNTO 124);
	wire_altbarrel_shift6_w_sbit_w_range281w <= sbit_w(30 DOWNTO 0);
	wire_altbarrel_shift6_w_sbit_w_range304w <= sbit_w(61 DOWNTO 31);
	wire_altbarrel_shift6_w_sbit_w_range324w <= sbit_w(92 DOWNTO 62);
	wire_altbarrel_shift6_w_sel_w_range286w(0) <= sel_w(0);
	wire_altbarrel_shift6_w_sel_w_range307w(0) <= sel_w(1);
	wire_altbarrel_shift6_w_sel_w_range329w(0) <= sel_w(2);
	wire_altbarrel_shift6_w_sel_w_range352w(0) <= sel_w(3);
	wire_altbarrel_shift6_w_sel_w_range371w(0) <= sel_w(4);
	wire_altbarrel_shift6_w_smux_w_range374w <= smux_w(154 DOWNTO 124);
	wire_altbarrel_shift6_w_smux_w_range333w <= smux_w(92 DOWNTO 62);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(4) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift6_w_smux_w_range333w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift6_w_smux_w_range374w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --converter_altbarrel_shift_svf

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 4 reg 185 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  converter_altfp_convert_tum IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (8 DOWNTO 0)
	 ); 
 END converter_altfp_convert_tum;

 ARCHITECTURE RTL OF converter_altfp_convert_tum IS

	 SIGNAL  wire_altbarrel_shift6_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL	 added_power2_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit1_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 below_lower_limit2_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit2_reg3_w_lg_q228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 below_lower_limit2_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_below_lower_limit2_reg4_w_lg_q259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 equal_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_equal_upper_limit_reg3_w_lg_q219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exceed_upper_limit_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exceed_upper_limit_reg3_w_lg_q220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exceed_upper_limit_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_and_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_or_reg4_w_lg_q117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 int_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 int_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_int_or_reg3_w_lg_q218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 integer_result_reg	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 integer_rounded_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lowest_int_sel_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_lowest_int_sel_reg_w_lg_q256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_or1_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or2_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_or_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_or_reg4_w_lg_q119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 mantissa_input_reg	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_exceeder_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 power2_value_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_input_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_input_reg3_w_lg_q221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sign_input_reg3_w_lg_q223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_input_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub7_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_w_lg_cout232w233w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_cout231w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub8_w_lg_cout232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub8_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub9_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr1_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_alb	:	STD_LOGIC;
	 SIGNAL  wire_max_shift_compare_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w200w201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_add_1_w205w206w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_below_limit_exceeders266w267w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exceed_limit_exceeders277w278w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w200w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_lowest_integer_selector212w213w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w237w270w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_input_w237w238w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w204w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders265w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders276w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector211w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w269w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w236w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range8w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range13w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range18w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range23w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range28w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range33w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_and_range38w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_add_1_w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_below_limit_exceeders266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_denormal_input_w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exceed_limit_exceeders277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_lowest_integer_selector212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_input_w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_input_w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_input_w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinity_input_w273w274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinity_input_w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range6w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range11w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range16w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range21w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range26w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range31w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_or_range36w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range47w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range74w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range71w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range68w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range65w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range62w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range59w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range56w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range53w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or1_range50w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range84w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range81w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range111w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range108w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range105w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range102w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range99w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range96w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range93w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range90w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_or2_range87w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range134w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range164w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range167w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range170w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range173w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range176w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range179w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range182w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range185w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range188w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range191w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range137w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range194w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range140w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range143w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range146w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range149w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range152w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range155w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range158w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_or_range161w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_cout_w :	STD_LOGIC;
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  all_zeroes_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  barrel_mantissa_input :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  barrel_zero_padding_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  below_limit_exceeders :	STD_LOGIC;
	 SIGNAL  below_limit_integer :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  below_lower_limit1_w :	STD_LOGIC;
	 SIGNAL  below_lower_limit2_w :	STD_LOGIC;
	 SIGNAL  bias_value_less_1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  denormal_input_w :	STD_LOGIC;
	 SIGNAL  equal_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exceed_limit_exceeders :	STD_LOGIC;
	 SIGNAL  exceed_limit_integer :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exceed_upper_limit_w :	STD_LOGIC;
	 SIGNAL  exp_and :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_and_w :	STD_LOGIC;
	 SIGNAL  exp_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or_w :	STD_LOGIC;
	 SIGNAL  exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  implied_mantissa_input :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  infinity_input_w :	STD_LOGIC;
	 SIGNAL  infinity_value_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  int_or1_w :	STD_LOGIC;
	 SIGNAL  integer_output :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  integer_post_round :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  integer_pre_round :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  integer_result :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  integer_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  integer_rounded_tmp :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  integer_tmp_output :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  inv_add_1_adder1_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  inv_add_1_adder2_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  inv_integer :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  lbarrel_shift_result_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  lbarrel_shift_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  lower_limit_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_selector :	STD_LOGIC;
	 SIGNAL  lowest_integer_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  man_bus1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_bus2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or1 :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  man_or1_w :	STD_LOGIC;
	 SIGNAL  man_or2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  man_or2_w :	STD_LOGIC;
	 SIGNAL  man_or_w :	STD_LOGIC;
	 SIGNAL  mantissa_input :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  max_shift_reg_w :	STD_LOGIC;
	 SIGNAL  max_shift_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  more_than_max_shift_w :	STD_LOGIC;
	 SIGNAL  nan_input_w :	STD_LOGIC;
	 SIGNAL  neg_infi_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  padded_exponent_input :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  pos_infi_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  power2_value_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  sign_input :	STD_LOGIC;
	 SIGNAL  sign_input_w :	STD_LOGIC;
	 SIGNAL  signed_integer :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  sticky_bus :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  sticky_or :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  unsigned_integer :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  upper_limit_w :	STD_LOGIC;
	 SIGNAL  zero_input_w :	STD_LOGIC;
	 SIGNAL  wire_w_exp_and_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_and_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bus_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_or_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_inv_integer_range217w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus1_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_bus2_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or1_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_or2_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bus_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_or_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  converter_altbarrel_shift_svf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w200w201w202w(0) <= wire_w_lg_w_lg_guard_bit_w200w201w(0) AND sticky_bit_w;
	loop25 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_add_1_w205w206w(i) <= wire_w_lg_add_1_w205w(0) AND integer_pre_round(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_below_limit_exceeders266w267w(i) <= wire_w_lg_below_limit_exceeders266w(0) AND integer_output(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_exceed_limit_exceeders277w278w(i) <= wire_w_lg_exceed_limit_exceeders277w(0) AND below_limit_integer(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_guard_bit_w200w201w(0) <= wire_w_lg_guard_bit_w200w(0) AND round_bit_w;
	loop28 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_lowest_integer_selector212w213w(i) <= wire_w_lg_lowest_integer_selector212w(0) AND integer_rounded_tmp(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_sign_input_w237w270w(i) <= wire_w_lg_sign_input_w237w(0) AND pos_infi_w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_sign_input_w237w238w(i) <= wire_w_lg_sign_input_w237w(0) AND unsigned_integer(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_add_1_w204w(i) <= add_1_w AND integer_post_round(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_below_limit_exceeders265w(i) <= below_limit_exceeders AND all_zeroes_w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_exceed_limit_exceeders276w(i) <= exceed_limit_exceeders AND infinity_value_w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_lowest_integer_selector211w(i) <= lowest_integer_selector AND lowest_integer_value(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_sign_input_w269w(i) <= sign_input_w AND neg_infi_w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_sign_input_w236w(i) <= sign_input_w AND signed_integer(i);
	END GENERATE loop36;
	wire_w_lg_w_exp_and_range8w14w(0) <= wire_w_exp_and_range8w(0) AND wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_and_range13w19w(0) <= wire_w_exp_and_range13w(0) AND wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_and_range18w24w(0) <= wire_w_exp_and_range18w(0) AND wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_and_range23w29w(0) <= wire_w_exp_and_range23w(0) AND wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_and_range28w34w(0) <= wire_w_exp_and_range28w(0) AND wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_and_range33w39w(0) <= wire_w_exp_and_range33w(0) AND wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_and_range38w44w(0) <= wire_w_exp_and_range38w(0) AND wire_w_exp_bus_range40w(0);
	wire_w_lg_add_1_w205w(0) <= NOT add_1_w;
	wire_w_lg_below_limit_exceeders266w(0) <= NOT below_limit_exceeders;
	wire_w_lg_denormal_input_w257w(0) <= NOT denormal_input_w;
	wire_w_lg_exceed_limit_exceeders277w(0) <= NOT exceed_limit_exceeders;
	wire_w_lg_guard_bit_w200w(0) <= NOT guard_bit_w;
	wire_w_lg_lowest_integer_selector212w(0) <= NOT lowest_integer_selector;
	wire_w_lg_nan_input_w272w(0) <= NOT nan_input_w;
	wire_w_lg_sign_input_w237w(0) <= NOT sign_input_w;
	wire_w_lg_zero_input_w258w(0) <= NOT zero_input_w;
	wire_w_lg_w_lg_infinity_input_w273w274w(0) <= wire_w_lg_infinity_input_w273w(0) OR exceed_upper_limit_reg4;
	wire_w_lg_infinity_input_w273w(0) <= infinity_input_w OR max_shift_exceeder_reg;
	wire_w_lg_w_exp_or_range6w12w(0) <= wire_w_exp_or_range6w(0) OR wire_w_exp_bus_range10w(0);
	wire_w_lg_w_exp_or_range11w17w(0) <= wire_w_exp_or_range11w(0) OR wire_w_exp_bus_range15w(0);
	wire_w_lg_w_exp_or_range16w22w(0) <= wire_w_exp_or_range16w(0) OR wire_w_exp_bus_range20w(0);
	wire_w_lg_w_exp_or_range21w27w(0) <= wire_w_exp_or_range21w(0) OR wire_w_exp_bus_range25w(0);
	wire_w_lg_w_exp_or_range26w32w(0) <= wire_w_exp_or_range26w(0) OR wire_w_exp_bus_range30w(0);
	wire_w_lg_w_exp_or_range31w37w(0) <= wire_w_exp_or_range31w(0) OR wire_w_exp_bus_range35w(0);
	wire_w_lg_w_exp_or_range36w42w(0) <= wire_w_exp_or_range36w(0) OR wire_w_exp_bus_range40w(0);
	wire_w_lg_w_man_or1_range47w51w(0) <= wire_w_man_or1_range47w(0) OR wire_w_man_bus1_range49w(0);
	wire_w_lg_w_man_or1_range74w78w(0) <= wire_w_man_or1_range74w(0) OR wire_w_man_bus1_range76w(0);
	wire_w_lg_w_man_or1_range71w75w(0) <= wire_w_man_or1_range71w(0) OR wire_w_man_bus1_range73w(0);
	wire_w_lg_w_man_or1_range68w72w(0) <= wire_w_man_or1_range68w(0) OR wire_w_man_bus1_range70w(0);
	wire_w_lg_w_man_or1_range65w69w(0) <= wire_w_man_or1_range65w(0) OR wire_w_man_bus1_range67w(0);
	wire_w_lg_w_man_or1_range62w66w(0) <= wire_w_man_or1_range62w(0) OR wire_w_man_bus1_range64w(0);
	wire_w_lg_w_man_or1_range59w63w(0) <= wire_w_man_or1_range59w(0) OR wire_w_man_bus1_range61w(0);
	wire_w_lg_w_man_or1_range56w60w(0) <= wire_w_man_or1_range56w(0) OR wire_w_man_bus1_range58w(0);
	wire_w_lg_w_man_or1_range53w57w(0) <= wire_w_man_or1_range53w(0) OR wire_w_man_bus1_range55w(0);
	wire_w_lg_w_man_or1_range50w54w(0) <= wire_w_man_or1_range50w(0) OR wire_w_man_bus1_range52w(0);
	wire_w_lg_w_man_or2_range84w88w(0) <= wire_w_man_or2_range84w(0) OR wire_w_man_bus2_range86w(0);
	wire_w_lg_w_man_or2_range81w85w(0) <= wire_w_man_or2_range81w(0) OR wire_w_man_bus2_range83w(0);
	wire_w_lg_w_man_or2_range111w115w(0) <= wire_w_man_or2_range111w(0) OR wire_w_man_bus2_range113w(0);
	wire_w_lg_w_man_or2_range108w112w(0) <= wire_w_man_or2_range108w(0) OR wire_w_man_bus2_range110w(0);
	wire_w_lg_w_man_or2_range105w109w(0) <= wire_w_man_or2_range105w(0) OR wire_w_man_bus2_range107w(0);
	wire_w_lg_w_man_or2_range102w106w(0) <= wire_w_man_or2_range102w(0) OR wire_w_man_bus2_range104w(0);
	wire_w_lg_w_man_or2_range99w103w(0) <= wire_w_man_or2_range99w(0) OR wire_w_man_bus2_range101w(0);
	wire_w_lg_w_man_or2_range96w100w(0) <= wire_w_man_or2_range96w(0) OR wire_w_man_bus2_range98w(0);
	wire_w_lg_w_man_or2_range93w97w(0) <= wire_w_man_or2_range93w(0) OR wire_w_man_bus2_range95w(0);
	wire_w_lg_w_man_or2_range90w94w(0) <= wire_w_man_or2_range90w(0) OR wire_w_man_bus2_range92w(0);
	wire_w_lg_w_man_or2_range87w91w(0) <= wire_w_man_or2_range87w(0) OR wire_w_man_bus2_range89w(0);
	wire_w_lg_w_sticky_or_range134w138w(0) <= wire_w_sticky_or_range134w(0) OR wire_w_sticky_bus_range136w(0);
	wire_w_lg_w_sticky_or_range164w168w(0) <= wire_w_sticky_or_range164w(0) OR wire_w_sticky_bus_range166w(0);
	wire_w_lg_w_sticky_or_range167w171w(0) <= wire_w_sticky_or_range167w(0) OR wire_w_sticky_bus_range169w(0);
	wire_w_lg_w_sticky_or_range170w174w(0) <= wire_w_sticky_or_range170w(0) OR wire_w_sticky_bus_range172w(0);
	wire_w_lg_w_sticky_or_range173w177w(0) <= wire_w_sticky_or_range173w(0) OR wire_w_sticky_bus_range175w(0);
	wire_w_lg_w_sticky_or_range176w180w(0) <= wire_w_sticky_or_range176w(0) OR wire_w_sticky_bus_range178w(0);
	wire_w_lg_w_sticky_or_range179w183w(0) <= wire_w_sticky_or_range179w(0) OR wire_w_sticky_bus_range181w(0);
	wire_w_lg_w_sticky_or_range182w186w(0) <= wire_w_sticky_or_range182w(0) OR wire_w_sticky_bus_range184w(0);
	wire_w_lg_w_sticky_or_range185w189w(0) <= wire_w_sticky_or_range185w(0) OR wire_w_sticky_bus_range187w(0);
	wire_w_lg_w_sticky_or_range188w192w(0) <= wire_w_sticky_or_range188w(0) OR wire_w_sticky_bus_range190w(0);
	wire_w_lg_w_sticky_or_range191w195w(0) <= wire_w_sticky_or_range191w(0) OR wire_w_sticky_bus_range193w(0);
	wire_w_lg_w_sticky_or_range137w141w(0) <= wire_w_sticky_or_range137w(0) OR wire_w_sticky_bus_range139w(0);
	wire_w_lg_w_sticky_or_range194w198w(0) <= wire_w_sticky_or_range194w(0) OR wire_w_sticky_bus_range196w(0);
	wire_w_lg_w_sticky_or_range140w144w(0) <= wire_w_sticky_or_range140w(0) OR wire_w_sticky_bus_range142w(0);
	wire_w_lg_w_sticky_or_range143w147w(0) <= wire_w_sticky_or_range143w(0) OR wire_w_sticky_bus_range145w(0);
	wire_w_lg_w_sticky_or_range146w150w(0) <= wire_w_sticky_or_range146w(0) OR wire_w_sticky_bus_range148w(0);
	wire_w_lg_w_sticky_or_range149w153w(0) <= wire_w_sticky_or_range149w(0) OR wire_w_sticky_bus_range151w(0);
	wire_w_lg_w_sticky_or_range152w156w(0) <= wire_w_sticky_or_range152w(0) OR wire_w_sticky_bus_range154w(0);
	wire_w_lg_w_sticky_or_range155w159w(0) <= wire_w_sticky_or_range155w(0) OR wire_w_sticky_bus_range157w(0);
	wire_w_lg_w_sticky_or_range158w162w(0) <= wire_w_sticky_or_range158w(0) OR wire_w_sticky_bus_range160w(0);
	wire_w_lg_w_sticky_or_range161w165w(0) <= wire_w_sticky_or_range161w(0) OR wire_w_sticky_bus_range163w(0);
	aclr <= '0';
	add_1_cout_w <= ((wire_add_sub7_cout AND add_1_w) AND wire_sign_input_reg3_w_lg_q223w(0));
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w200w201w202w(0) OR (guard_bit_w AND round_bit_w));
	all_zeroes_w <= ( "0" & "00000000");
	barrel_mantissa_input <= ( barrel_zero_padding_w & implied_mantissa_input);
	barrel_zero_padding_w <= (OTHERS => '0');
	below_limit_exceeders <= (((denormal_input_w OR zero_input_w) OR lower_limit_selector) OR nan_input_w);
	below_limit_integer <= (wire_w_lg_w_lg_below_limit_exceeders266w267w OR wire_w_lg_below_limit_exceeders265w);
	below_lower_limit1_w <= wire_cmpr2_aeb;
	below_lower_limit2_w <= wire_cmpr3_alb;
	bias_value_less_1_w <= "01111110";
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_res_w <= "10000111";
	denormal_input_w <= (wire_exp_or_reg4_w_lg_q117w(0) AND man_or_reg4);
	equal_upper_limit_w <= wire_cmpr1_aeb;
	exceed_limit_exceeders <= (wire_w_lg_w_lg_infinity_input_w273w274w(0) AND wire_w_lg_nan_input_w272w(0));
	exceed_limit_integer <= (wire_w_lg_w_lg_exceed_limit_exceeders277w278w OR wire_w_lg_exceed_limit_exceeders276w);
	exceed_upper_limit_w <= wire_cmpr1_agb;
	exp_and <= ( wire_w_lg_w_exp_and_range38w44w & wire_w_lg_w_exp_and_range33w39w & wire_w_lg_w_exp_and_range28w34w & wire_w_lg_w_exp_and_range23w29w & wire_w_lg_w_exp_and_range18w24w & wire_w_lg_w_exp_and_range13w19w & wire_w_lg_w_exp_and_range8w14w & exp_bus(0));
	exp_and_w <= exp_and(7);
	exp_bus <= exponent_input;
	exp_or <= ( wire_w_lg_w_exp_or_range36w42w & wire_w_lg_w_exp_or_range31w37w & wire_w_lg_w_exp_or_range26w32w & wire_w_lg_w_exp_or_range21w27w & wire_w_lg_w_exp_or_range16w22w & wire_w_lg_w_exp_or_range11w17w & wire_w_lg_w_exp_or_range6w12w & exp_bus(0));
	exp_or_w <= exp_or(7);
	exponent_input <= dataa_reg(30 DOWNTO 23);
	guard_bit_w <= wire_altbarrel_shift6_result(23);
	implied_mantissa_input <= ( "1" & mantissa_input_reg);
	infinity_input_w <= (exp_and_reg4 AND wire_man_or_reg4_w_lg_q119w(0));
	infinity_value_w <= (wire_w_lg_w_lg_sign_input_w237w270w OR wire_w_lg_sign_input_w269w);
	int_or1_w <= man_or2(4);
	integer_output <= ( sign_input_w & integer_tmp_output);
	integer_post_round <= wire_add_sub7_result;
	integer_pre_round <= lbarrel_shift_w;
	integer_result <= exceed_limit_integer;
	integer_rounded <= (wire_w_lg_w_lg_lowest_integer_selector212w213w OR wire_w_lg_lowest_integer_selector211w);
	integer_rounded_tmp <= (wire_w_lg_w_lg_add_1_w205w206w OR wire_w_lg_add_1_w204w);
	integer_tmp_output <= (wire_w_lg_w_lg_sign_input_w237w238w OR wire_w_lg_sign_input_w236w);
	inv_add_1_adder1_w <= wire_add_sub8_result;
	inv_add_1_adder2_w <= (wire_add_sub8_w_lg_w_lg_cout232w233w OR wire_add_sub8_w_lg_cout231w);
	inv_integer <= (NOT integer_rounded_reg);
	lbarrel_shift_result_w <= wire_altbarrel_shift6_result;
	lbarrel_shift_w <= lbarrel_shift_result_w(30 DOWNTO 23);
	lower_limit_selector <= ((wire_below_lower_limit2_reg4_w_lg_q259w(0) AND wire_w_lg_denormal_input_w257w(0)) AND wire_lowest_int_sel_reg_w_lg_q256w(0));
	lowest_integer_selector <= (below_lower_limit1_reg3 AND man_or_reg3);
	lowest_integer_value <= ( barrel_zero_padding_w & "1");
	man_bus1 <= mantissa_input(10 DOWNTO 0);
	man_bus2 <= mantissa_input(22 DOWNTO 11);
	man_or1 <= ( man_bus1(10) & wire_w_lg_w_man_or1_range47w51w & wire_w_lg_w_man_or1_range50w54w & wire_w_lg_w_man_or1_range53w57w & wire_w_lg_w_man_or1_range56w60w & wire_w_lg_w_man_or1_range59w63w & wire_w_lg_w_man_or1_range62w66w & wire_w_lg_w_man_or1_range65w69w & wire_w_lg_w_man_or1_range68w72w & wire_w_lg_w_man_or1_range71w75w & wire_w_lg_w_man_or1_range74w78w);
	man_or1_w <= man_or1(0);
	man_or2 <= ( man_bus2(11) & wire_w_lg_w_man_or2_range81w85w & wire_w_lg_w_man_or2_range84w88w & wire_w_lg_w_man_or2_range87w91w & wire_w_lg_w_man_or2_range90w94w & wire_w_lg_w_man_or2_range93w97w & wire_w_lg_w_man_or2_range96w100w & wire_w_lg_w_man_or2_range99w103w & wire_w_lg_w_man_or2_range102w106w & wire_w_lg_w_man_or2_range105w109w & wire_w_lg_w_man_or2_range108w112w & wire_w_lg_w_man_or2_range111w115w);
	man_or2_w <= man_or2(0);
	man_or_w <= (man_or1_reg1 OR man_or2_reg1);
	mantissa_input <= dataa_reg(22 DOWNTO 0);
	max_shift_reg_w <= max_shift_reg;
	max_shift_w <= "00111";
	more_than_max_shift_w <= ((max_shift_reg_w AND add_1_cout_w) AND wire_below_lower_limit2_reg3_w_lg_q228w(0));
	nan_input_w <= (exp_and_reg4 AND man_or_reg4);
	neg_infi_w <= ( "1" & "00000000");
	padded_exponent_input <= exponent_input;
	pos_infi_w <= ( "0" & "11111111");
	power2_value_w <= wire_add_sub4_result(4 DOWNTO 0);
	result <= result_w;
	result_w <= integer_result_reg;
	round_bit_w <= wire_altbarrel_shift6_result(22);
	sign_input <= dataa_reg(31);
	sign_input_w <= sign_input_reg4;
	signed_integer <= ( inv_add_1_adder2_w & inv_add_1_adder1_w);
	sticky_bit_w <= sticky_or(21);
	sticky_bus <= wire_altbarrel_shift6_result(21 DOWNTO 0);
	sticky_or <= ( wire_w_lg_w_sticky_or_range194w198w & wire_w_lg_w_sticky_or_range191w195w & wire_w_lg_w_sticky_or_range188w192w & wire_w_lg_w_sticky_or_range185w189w & wire_w_lg_w_sticky_or_range182w186w & wire_w_lg_w_sticky_or_range179w183w & wire_w_lg_w_sticky_or_range176w180w & wire_w_lg_w_sticky_or_range173w177w & wire_w_lg_w_sticky_or_range170w174w & wire_w_lg_w_sticky_or_range167w171w & wire_w_lg_w_sticky_or_range164w168w & wire_w_lg_w_sticky_or_range161w165w & wire_w_lg_w_sticky_or_range158w162w & wire_w_lg_w_sticky_or_range155w159w & wire_w_lg_w_sticky_or_range152w156w & wire_w_lg_w_sticky_or_range149w153w & wire_w_lg_w_sticky_or_range146w150w & wire_w_lg_w_sticky_or_range143w147w & wire_w_lg_w_sticky_or_range140w144w & wire_w_lg_w_sticky_or_range137w141w & wire_w_lg_w_sticky_or_range134w138w & sticky_bus(0));
	unsigned_integer <= integer_rounded_reg;
	upper_limit_w <= ((wire_sign_input_reg3_w_lg_q223w(0) AND (exceed_upper_limit_reg3 OR equal_upper_limit_reg3)) OR wire_sign_input_reg3_w_lg_q221w(0));
	zero_input_w <= (wire_exp_or_reg4_w_lg_q117w(0) AND wire_man_or_reg4_w_lg_q119w(0));
	wire_w_exp_and_range8w(0) <= exp_and(0);
	wire_w_exp_and_range13w(0) <= exp_and(1);
	wire_w_exp_and_range18w(0) <= exp_and(2);
	wire_w_exp_and_range23w(0) <= exp_and(3);
	wire_w_exp_and_range28w(0) <= exp_and(4);
	wire_w_exp_and_range33w(0) <= exp_and(5);
	wire_w_exp_and_range38w(0) <= exp_and(6);
	wire_w_exp_bus_range10w(0) <= exp_bus(1);
	wire_w_exp_bus_range15w(0) <= exp_bus(2);
	wire_w_exp_bus_range20w(0) <= exp_bus(3);
	wire_w_exp_bus_range25w(0) <= exp_bus(4);
	wire_w_exp_bus_range30w(0) <= exp_bus(5);
	wire_w_exp_bus_range35w(0) <= exp_bus(6);
	wire_w_exp_bus_range40w(0) <= exp_bus(7);
	wire_w_exp_or_range6w(0) <= exp_or(0);
	wire_w_exp_or_range11w(0) <= exp_or(1);
	wire_w_exp_or_range16w(0) <= exp_or(2);
	wire_w_exp_or_range21w(0) <= exp_or(3);
	wire_w_exp_or_range26w(0) <= exp_or(4);
	wire_w_exp_or_range31w(0) <= exp_or(5);
	wire_w_exp_or_range36w(0) <= exp_or(6);
	wire_w_inv_integer_range217w <= inv_integer(7 DOWNTO 4);
	wire_w_man_bus1_range76w(0) <= man_bus1(0);
	wire_w_man_bus1_range73w(0) <= man_bus1(1);
	wire_w_man_bus1_range70w(0) <= man_bus1(2);
	wire_w_man_bus1_range67w(0) <= man_bus1(3);
	wire_w_man_bus1_range64w(0) <= man_bus1(4);
	wire_w_man_bus1_range61w(0) <= man_bus1(5);
	wire_w_man_bus1_range58w(0) <= man_bus1(6);
	wire_w_man_bus1_range55w(0) <= man_bus1(7);
	wire_w_man_bus1_range52w(0) <= man_bus1(8);
	wire_w_man_bus1_range49w(0) <= man_bus1(9);
	wire_w_man_bus2_range113w(0) <= man_bus2(0);
	wire_w_man_bus2_range83w(0) <= man_bus2(10);
	wire_w_man_bus2_range110w(0) <= man_bus2(1);
	wire_w_man_bus2_range107w(0) <= man_bus2(2);
	wire_w_man_bus2_range104w(0) <= man_bus2(3);
	wire_w_man_bus2_range101w(0) <= man_bus2(4);
	wire_w_man_bus2_range98w(0) <= man_bus2(5);
	wire_w_man_bus2_range95w(0) <= man_bus2(6);
	wire_w_man_bus2_range92w(0) <= man_bus2(7);
	wire_w_man_bus2_range89w(0) <= man_bus2(8);
	wire_w_man_bus2_range86w(0) <= man_bus2(9);
	wire_w_man_or1_range47w(0) <= man_or1(10);
	wire_w_man_or1_range74w(0) <= man_or1(1);
	wire_w_man_or1_range71w(0) <= man_or1(2);
	wire_w_man_or1_range68w(0) <= man_or1(3);
	wire_w_man_or1_range65w(0) <= man_or1(4);
	wire_w_man_or1_range62w(0) <= man_or1(5);
	wire_w_man_or1_range59w(0) <= man_or1(6);
	wire_w_man_or1_range56w(0) <= man_or1(7);
	wire_w_man_or1_range53w(0) <= man_or1(8);
	wire_w_man_or1_range50w(0) <= man_or1(9);
	wire_w_man_or2_range84w(0) <= man_or2(10);
	wire_w_man_or2_range81w(0) <= man_or2(11);
	wire_w_man_or2_range111w(0) <= man_or2(1);
	wire_w_man_or2_range108w(0) <= man_or2(2);
	wire_w_man_or2_range105w(0) <= man_or2(3);
	wire_w_man_or2_range102w(0) <= man_or2(4);
	wire_w_man_or2_range99w(0) <= man_or2(5);
	wire_w_man_or2_range96w(0) <= man_or2(6);
	wire_w_man_or2_range93w(0) <= man_or2(7);
	wire_w_man_or2_range90w(0) <= man_or2(8);
	wire_w_man_or2_range87w(0) <= man_or2(9);
	wire_w_sticky_bus_range163w(0) <= sticky_bus(10);
	wire_w_sticky_bus_range166w(0) <= sticky_bus(11);
	wire_w_sticky_bus_range169w(0) <= sticky_bus(12);
	wire_w_sticky_bus_range172w(0) <= sticky_bus(13);
	wire_w_sticky_bus_range175w(0) <= sticky_bus(14);
	wire_w_sticky_bus_range178w(0) <= sticky_bus(15);
	wire_w_sticky_bus_range181w(0) <= sticky_bus(16);
	wire_w_sticky_bus_range184w(0) <= sticky_bus(17);
	wire_w_sticky_bus_range187w(0) <= sticky_bus(18);
	wire_w_sticky_bus_range190w(0) <= sticky_bus(19);
	wire_w_sticky_bus_range136w(0) <= sticky_bus(1);
	wire_w_sticky_bus_range193w(0) <= sticky_bus(20);
	wire_w_sticky_bus_range196w(0) <= sticky_bus(21);
	wire_w_sticky_bus_range139w(0) <= sticky_bus(2);
	wire_w_sticky_bus_range142w(0) <= sticky_bus(3);
	wire_w_sticky_bus_range145w(0) <= sticky_bus(4);
	wire_w_sticky_bus_range148w(0) <= sticky_bus(5);
	wire_w_sticky_bus_range151w(0) <= sticky_bus(6);
	wire_w_sticky_bus_range154w(0) <= sticky_bus(7);
	wire_w_sticky_bus_range157w(0) <= sticky_bus(8);
	wire_w_sticky_bus_range160w(0) <= sticky_bus(9);
	wire_w_sticky_or_range134w(0) <= sticky_or(0);
	wire_w_sticky_or_range164w(0) <= sticky_or(10);
	wire_w_sticky_or_range167w(0) <= sticky_or(11);
	wire_w_sticky_or_range170w(0) <= sticky_or(12);
	wire_w_sticky_or_range173w(0) <= sticky_or(13);
	wire_w_sticky_or_range176w(0) <= sticky_or(14);
	wire_w_sticky_or_range179w(0) <= sticky_or(15);
	wire_w_sticky_or_range182w(0) <= sticky_or(16);
	wire_w_sticky_or_range185w(0) <= sticky_or(17);
	wire_w_sticky_or_range188w(0) <= sticky_or(18);
	wire_w_sticky_or_range191w(0) <= sticky_or(19);
	wire_w_sticky_or_range137w(0) <= sticky_or(1);
	wire_w_sticky_or_range194w(0) <= sticky_or(20);
	wire_w_sticky_or_range140w(0) <= sticky_or(2);
	wire_w_sticky_or_range143w(0) <= sticky_or(3);
	wire_w_sticky_or_range146w(0) <= sticky_or(4);
	wire_w_sticky_or_range149w(0) <= sticky_or(5);
	wire_w_sticky_or_range152w(0) <= sticky_or(6);
	wire_w_sticky_or_range155w(0) <= sticky_or(7);
	wire_w_sticky_or_range158w(0) <= sticky_or(8);
	wire_w_sticky_or_range161w(0) <= sticky_or(9);
	altbarrel_shift6 :  converter_altbarrel_shift_svf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => barrel_mantissa_input,
		distance => power2_value_reg,
		result => wire_altbarrel_shift6_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN added_power2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN added_power2_reg <= wire_add_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg1 <= below_lower_limit1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg2 <= below_lower_limit1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit1_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit1_reg3 <= below_lower_limit1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg1 <= below_lower_limit2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg2 <= below_lower_limit2_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg3 <= below_lower_limit2_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit2_reg3_w_lg_q228w(0) <= NOT below_lower_limit2_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN below_lower_limit2_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN below_lower_limit2_reg4 <= below_lower_limit2_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_below_lower_limit2_reg4_w_lg_q259w(0) <= below_lower_limit2_reg4 AND wire_w_lg_zero_input_w258w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_reg <= dataa;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg1 <= equal_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg2 <= equal_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN equal_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN equal_upper_limit_reg3 <= equal_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_equal_upper_limit_reg3_w_lg_q219w(0) <= equal_upper_limit_reg3 AND wire_int_or_reg3_w_lg_q218w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg1 <= exceed_upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg2 <= exceed_upper_limit_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg3 <= exceed_upper_limit_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_exceed_upper_limit_reg3_w_lg_q220w(0) <= exceed_upper_limit_reg3 OR wire_equal_upper_limit_reg3_w_lg_q219w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exceed_upper_limit_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exceed_upper_limit_reg4 <= upper_limit_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg1 <= exp_and_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg2 <= exp_and_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg3 <= exp_and_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_and_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_and_reg4 <= exp_and_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg1 <= exp_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg2 <= exp_or_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg3 <= exp_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_or_reg4 <= exp_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_or_reg4_w_lg_q117w(0) <= NOT exp_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or1_reg1 <= int_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg2 <= int_or1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN int_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN int_or_reg3 <= int_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_int_or_reg3_w_lg_q218w(0) <= int_or_reg3 OR add_1_w;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_result_reg <= integer_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN integer_rounded_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN integer_rounded_reg <= integer_rounded;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lowest_int_sel_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lowest_int_sel_reg <= lowest_integer_selector;
			END IF;
		END IF;
	END PROCESS;
	wire_lowest_int_sel_reg_w_lg_q256w(0) <= NOT lowest_int_sel_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or1_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or1_reg1 <= man_or1_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or2_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or2_reg1 <= man_or2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg2 <= man_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg3 <= man_or_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_or_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_or_reg4 <= man_or_reg3;
			END IF;
		END IF;
	END PROCESS;
	wire_man_or_reg4_w_lg_q119w(0) <= NOT man_or_reg4;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_input_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_input_reg <= mantissa_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_exceeder_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_exceeder_reg <= more_than_max_shift_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN max_shift_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN max_shift_reg <= wire_max_shift_compare_agb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN power2_value_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN power2_value_reg <= power2_value_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg1 <= sign_input;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg2 <= sign_input_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg3 <= sign_input_reg2;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_input_reg3_w_lg_q221w(0) <= sign_input_reg3 AND wire_exceed_upper_limit_reg3_w_lg_q220w(0);
	wire_sign_input_reg3_w_lg_q223w(0) <= NOT sign_input_reg3;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_input_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_input_reg4 <= sign_input_reg3;
			END IF;
		END IF;
	END PROCESS;
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_input,
		datab => bias_value_w,
		result => wire_add_sub4_result
	  );
	wire_add_sub5_datab <= "00001";
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 5,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => power2_value_reg,
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub7_datab <= "00000001";
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub7_cout,
		dataa => integer_pre_round,
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_add_sub8_w_lg_w_lg_cout232w233w(i) <= wire_add_sub8_w_lg_cout232w(0) AND wire_w_inv_integer_range217w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_add_sub8_w_lg_cout231w(i) <= wire_add_sub8_cout AND wire_add_sub9_result(i);
	END GENERATE loop38;
	wire_add_sub8_w_lg_cout232w(0) <= NOT wire_add_sub8_cout;
	wire_add_sub8_datab <= "0001";
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 4,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub8_cout,
		dataa => inv_integer(3 DOWNTO 0),
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	wire_add_sub9_datab <= "0001";
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 4,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => inv_integer(7 DOWNTO 4),
		datab => wire_add_sub9_datab,
		result => wire_add_sub9_result
	  );
	cmpr1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr1_aeb,
		agb => wire_cmpr1_agb,
		dataa => padded_exponent_input,
		datab => const_bias_value_add_width_res_w
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr2_aeb,
		dataa => exponent_input,
		datab => bias_value_less_1_w
	  );
	cmpr3 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr3_alb,
		dataa => exponent_input,
		datab => bias_value_w
	  );
	max_shift_compare :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		agb => wire_max_shift_compare_agb,
		dataa => added_power2_reg,
		datab => max_shift_w
	  );

 END RTL; --converter_altfp_convert_tum
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY converter IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0)
	);
END converter;


ARCHITECTURE RTL OF converter IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (8 DOWNTO 0);



	COMPONENT converter_altfp_convert_tum
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (8 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(8 DOWNTO 0);

	converter_altfp_convert_tum_component : converter_altfp_convert_tum
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "FLOAT2INT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "9"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "9"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 9 0 OUTPUT NODEFVAL "result[8..0]"
-- Retrieval info: CONNECT: result 0 0 9 0 @result 0 0 9 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL converter.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: lpm
